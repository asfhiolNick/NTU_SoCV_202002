// RTL (Verilog) generated @ Mon Mar  8 04:38:47 2021 by V3 
//               compiled @ Mar  8 2021 00:47:13
// Internal nets are renamed with prefix "v3_1615207127_".

// Module vendingMachine
module vendingMachine
(
   clk,
   reset,
   coinInA,
   coinInB,
   coinInC,
   coinInD,
   itemTypeIn,
   itemNumberIn,
   forceIn,
   coinOutA,
   coinOutB,
   coinOutC,
   coinOutD,
   itemTypeOut,
   itemNumberOut,
   serviceTypeOut
);

   // Clock Signal for Synchronous DFF
   input clk;

   // I/O Declarations
   input reset;
   input [5:0] coinInA;
   input [5:0] coinInB;
   input [5:0] coinInC;
   input [5:0] coinInD;
   input [1:0] itemTypeIn;
   input [2:0] itemNumberIn;
   input forceIn;
   output [5:0] coinOutA;
   output [5:0] coinOutB;
   output [5:0] coinOutC;
   output [5:0] coinOutD;
   output [1:0] itemTypeOut;
   output [2:0] itemNumberOut;
   output [1:0] serviceTypeOut;

   // Wire and Reg Declarations
   wire v3_1615207127_0;
   wire clk;
   wire reset;
   wire [5:0] coinInA;
   wire [5:0] coinInB;
   wire [5:0] coinInC;
   wire [5:0] coinInD;
   wire [1:0] itemTypeIn;
   wire [2:0] itemNumberIn;
   wire forceIn;
   reg [5:0] v3_1615207127_10;
   reg [5:0] v3_1615207127_11;
   reg [5:0] v3_1615207127_12;
   reg [5:0] v3_1615207127_13;
   reg [1:0] v3_1615207127_14;
   reg [2:0] v3_1615207127_15;
   reg [1:0] v3_1615207127_16;
   reg v3_1615207127_17;
   reg v3_1615207127_18;
   reg [1:0] v3_1615207127_19;
   reg v3_1615207127_20;
   reg [12:0] v3_1615207127_21;
   reg [12:0] v3_1615207127_22;
   reg [5:0] v3_1615207127_23;
   reg [5:0] v3_1615207127_24;
   reg [5:0] v3_1615207127_25;
   reg [5:0] v3_1615207127_26;
   wire [5:0] v3_1615207127_27;
   wire [5:0] v3_1615207127_28;
   wire [5:0] v3_1615207127_29;
   wire [5:0] v3_1615207127_30;
   wire [5:0] v3_1615207127_31;
   wire [5:0] v3_1615207127_32;
   wire [5:0] v3_1615207127_33;
   wire [5:0] v3_1615207127_34;
   wire [5:0] v3_1615207127_35;
   wire [5:0] v3_1615207127_36;
   wire [5:0] v3_1615207127_37;
   wire [5:0] v3_1615207127_38;
   wire [5:0] v3_1615207127_39;
   wire [5:0] v3_1615207127_40;
   wire [5:0] v3_1615207127_41;
   wire v3_1615207127_42;
   wire v3_1615207127_43;
   wire [12:0] v3_1615207127_44;
   wire [5:0] v3_1615207127_45;
   wire v3_1615207127_46;
   wire [1:0] v3_1615207127_47;
   wire [5:0] v3_1615207127_48;
   wire v3_1615207127_49;
   wire [1:0] v3_1615207127_50;
   wire [5:0] v3_1615207127_51;
   wire [5:0] v3_1615207127_52;
   wire [5:0] v3_1615207127_53;
   wire [5:0] v3_1615207127_54;
   wire [5:0] v3_1615207127_55;
   wire [5:0] v3_1615207127_56;
   wire [5:0] v3_1615207127_57;
   wire v3_1615207127_58;
   wire v3_1615207127_59;
   wire [12:0] v3_1615207127_60;
   wire v3_1615207127_61;
   wire [1:0] v3_1615207127_62;
   wire [5:0] v3_1615207127_63;
   wire v3_1615207127_64;
   wire [5:0] v3_1615207127_65;
   wire v3_1615207127_66;
   wire [5:0] v3_1615207127_67;
   wire [5:0] v3_1615207127_68;
   wire [5:0] v3_1615207127_69;
   wire v3_1615207127_70;
   wire v3_1615207127_71;
   wire [2:0] v3_1615207127_72;
   wire v3_1615207127_73;
   wire [5:0] v3_1615207127_74;
   wire v3_1615207127_75;
   wire [5:0] v3_1615207127_76;
   wire [5:0] v3_1615207127_77;
   wire [5:0] v3_1615207127_78;
   wire [5:0] v3_1615207127_79;
   wire [5:0] v3_1615207127_80;
   wire [5:0] v3_1615207127_81;
   wire [5:0] v3_1615207127_82;
   wire [5:0] v3_1615207127_83;
   wire [5:0] v3_1615207127_84;
   wire [5:0] v3_1615207127_85;
   wire [5:0] v3_1615207127_86;
   wire [5:0] v3_1615207127_87;
   wire [5:0] v3_1615207127_88;
   wire [5:0] v3_1615207127_89;
   wire [5:0] v3_1615207127_90;
   wire [5:0] v3_1615207127_91;
   wire [5:0] v3_1615207127_92;
   wire [5:0] v3_1615207127_93;
   wire [5:0] v3_1615207127_94;
   wire [5:0] v3_1615207127_95;
   wire [5:0] v3_1615207127_96;
   wire [5:0] v3_1615207127_97;
   wire v3_1615207127_98;
   wire v3_1615207127_99;
   wire [12:0] v3_1615207127_100;
   wire [5:0] v3_1615207127_101;
   wire [5:0] v3_1615207127_102;
   wire [5:0] v3_1615207127_103;
   wire [5:0] v3_1615207127_104;
   wire [5:0] v3_1615207127_105;
   wire [5:0] v3_1615207127_106;
   wire [5:0] v3_1615207127_107;
   wire [5:0] v3_1615207127_108;
   wire [5:0] v3_1615207127_109;
   wire [5:0] v3_1615207127_110;
   wire [5:0] v3_1615207127_111;
   wire [5:0] v3_1615207127_112;
   wire [5:0] v3_1615207127_113;
   wire [5:0] v3_1615207127_114;
   wire [5:0] v3_1615207127_115;
   wire [5:0] v3_1615207127_116;
   wire [5:0] v3_1615207127_117;
   wire [5:0] v3_1615207127_118;
   wire [5:0] v3_1615207127_119;
   wire [5:0] v3_1615207127_120;
   wire [5:0] v3_1615207127_121;
   wire [5:0] v3_1615207127_122;
   wire [5:0] v3_1615207127_123;
   wire [5:0] v3_1615207127_124;
   wire [5:0] v3_1615207127_125;
   wire [5:0] v3_1615207127_126;
   wire [5:0] v3_1615207127_127;
   wire [5:0] v3_1615207127_128;
   wire v3_1615207127_129;
   wire v3_1615207127_130;
   wire [12:0] v3_1615207127_131;
   wire [5:0] v3_1615207127_132;
   wire [5:0] v3_1615207127_133;
   wire [5:0] v3_1615207127_134;
   wire [5:0] v3_1615207127_135;
   wire [5:0] v3_1615207127_136;
   wire [5:0] v3_1615207127_137;
   wire [5:0] v3_1615207127_138;
   wire [5:0] v3_1615207127_139;
   wire [5:0] v3_1615207127_140;
   wire [5:0] v3_1615207127_141;
   wire [5:0] v3_1615207127_142;
   wire [5:0] v3_1615207127_143;
   wire [5:0] v3_1615207127_144;
   wire [5:0] v3_1615207127_145;
   wire [5:0] v3_1615207127_146;
   wire [5:0] v3_1615207127_147;
   wire [5:0] v3_1615207127_148;
   wire [5:0] v3_1615207127_149;
   wire [5:0] v3_1615207127_150;
   wire [5:0] v3_1615207127_151;
   wire [5:0] v3_1615207127_152;
   wire [5:0] v3_1615207127_153;
   wire [5:0] v3_1615207127_154;
   wire [5:0] v3_1615207127_155;
   wire [5:0] v3_1615207127_156;
   wire [5:0] v3_1615207127_157;
   wire [5:0] v3_1615207127_158;
   wire [5:0] v3_1615207127_159;
   wire [5:0] v3_1615207127_160;
   wire [5:0] v3_1615207127_161;
   wire [5:0] v3_1615207127_162;
   wire [5:0] v3_1615207127_163;
   wire [5:0] v3_1615207127_164;
   wire [5:0] v3_1615207127_165;
   wire [1:0] v3_1615207127_166;
   wire [1:0] v3_1615207127_167;
   wire [1:0] v3_1615207127_168;
   wire [1:0] v3_1615207127_169;
   wire [1:0] v3_1615207127_170;
   wire [1:0] v3_1615207127_171;
   wire [1:0] v3_1615207127_172;
   wire [1:0] v3_1615207127_173;
   wire [1:0] v3_1615207127_174;
   wire [1:0] v3_1615207127_175;
   wire [2:0] v3_1615207127_176;
   wire [2:0] v3_1615207127_177;
   wire [2:0] v3_1615207127_178;
   wire [2:0] v3_1615207127_179;
   wire [2:0] v3_1615207127_180;
   wire [2:0] v3_1615207127_181;
   wire [2:0] v3_1615207127_182;
   wire [2:0] v3_1615207127_183;
   wire [2:0] v3_1615207127_184;
   wire [2:0] v3_1615207127_185;
   wire [2:0] v3_1615207127_186;
   wire [2:0] v3_1615207127_187;
   wire [2:0] v3_1615207127_188;
   wire [2:0] v3_1615207127_189;
   wire [2:0] v3_1615207127_190;
   wire [2:0] v3_1615207127_191;
   wire [2:0] v3_1615207127_192;
   wire [2:0] v3_1615207127_193;
   wire [2:0] v3_1615207127_194;
   wire [2:0] v3_1615207127_195;
   wire [2:0] v3_1615207127_196;
   wire [2:0] v3_1615207127_197;
   wire [2:0] v3_1615207127_198;
   wire [2:0] v3_1615207127_199;
   wire [2:0] v3_1615207127_200;
   wire v3_1615207127_201;
   wire v3_1615207127_202;
   wire [2:0] v3_1615207127_203;
   wire [2:0] v3_1615207127_204;
   wire [2:0] v3_1615207127_205;
   wire [2:0] v3_1615207127_206;
   wire [2:0] v3_1615207127_207;
   wire [2:0] v3_1615207127_208;
   wire [1:0] v3_1615207127_209;
   wire [1:0] v3_1615207127_210;
   wire [1:0] v3_1615207127_211;
   wire [1:0] v3_1615207127_212;
   wire [1:0] v3_1615207127_213;
   wire [1:0] v3_1615207127_214;
   wire [1:0] v3_1615207127_215;
   wire [1:0] v3_1615207127_216;
   wire [1:0] v3_1615207127_217;
   wire [1:0] v3_1615207127_218;
   wire [1:0] v3_1615207127_219;
   wire [1:0] v3_1615207127_220;
   wire [1:0] v3_1615207127_221;
   wire [1:0] v3_1615207127_222;
   wire [1:0] v3_1615207127_223;
   wire [1:0] v3_1615207127_224;
   wire [1:0] v3_1615207127_225;
   wire [1:0] v3_1615207127_226;
   wire [1:0] v3_1615207127_227;
   wire [1:0] v3_1615207127_228;
   wire [1:0] v3_1615207127_229;
   wire [1:0] v3_1615207127_230;
   wire v3_1615207127_231;
   wire v3_1615207127_232;
   wire v3_1615207127_233;
   wire v3_1615207127_234;
   wire v3_1615207127_235;
   wire v3_1615207127_236;
   wire v3_1615207127_237;
   wire v3_1615207127_238;
   wire v3_1615207127_239;
   wire v3_1615207127_240;
   wire v3_1615207127_241;
   wire v3_1615207127_242;
   wire v3_1615207127_243;
   wire v3_1615207127_244;
   wire v3_1615207127_245;
   wire v3_1615207127_246;
   wire v3_1615207127_247;
   wire v3_1615207127_248;
   wire v3_1615207127_249;
   wire v3_1615207127_250;
   wire v3_1615207127_251;
   wire v3_1615207127_252;
   wire v3_1615207127_253;
   wire v3_1615207127_254;
   wire [1:0] v3_1615207127_255;
   wire [1:0] v3_1615207127_256;
   wire [1:0] v3_1615207127_257;
   wire [1:0] v3_1615207127_258;
   wire [1:0] v3_1615207127_259;
   wire [1:0] v3_1615207127_260;
   wire [1:0] v3_1615207127_261;
   wire [1:0] v3_1615207127_262;
   wire [1:0] v3_1615207127_263;
   wire [1:0] v3_1615207127_264;
   wire [1:0] v3_1615207127_265;
   wire [1:0] v3_1615207127_266;
   wire [1:0] v3_1615207127_267;
   wire [1:0] v3_1615207127_268;
   wire [1:0] v3_1615207127_269;
   wire [1:0] v3_1615207127_270;
   wire [1:0] v3_1615207127_271;
   wire [1:0] v3_1615207127_272;
   wire [1:0] v3_1615207127_273;
   wire [1:0] v3_1615207127_274;
   wire [1:0] v3_1615207127_275;
   wire [1:0] v3_1615207127_276;
   wire [1:0] v3_1615207127_277;
   wire [1:0] v3_1615207127_278;
   wire [1:0] v3_1615207127_279;
   wire [1:0] v3_1615207127_280;
   wire [1:0] v3_1615207127_281;
   wire [1:0] v3_1615207127_282;
   wire [1:0] v3_1615207127_283;
   wire [1:0] v3_1615207127_284;
   wire [1:0] v3_1615207127_285;
   wire [1:0] v3_1615207127_286;
   wire [1:0] v3_1615207127_287;
   wire [1:0] v3_1615207127_288;
   wire [1:0] v3_1615207127_289;
   wire [1:0] v3_1615207127_290;
   wire [1:0] v3_1615207127_291;
   wire v3_1615207127_292;
   wire v3_1615207127_293;
   wire v3_1615207127_294;
   wire v3_1615207127_295;
   wire v3_1615207127_296;
   wire v3_1615207127_297;
   wire v3_1615207127_298;
   wire v3_1615207127_299;
   wire v3_1615207127_300;
   wire v3_1615207127_301;
   wire [12:0] v3_1615207127_302;
   wire [12:0] v3_1615207127_303;
   wire [12:0] v3_1615207127_304;
   wire [12:0] v3_1615207127_305;
   wire [12:0] v3_1615207127_306;
   wire [12:0] v3_1615207127_307;
   wire [12:0] v3_1615207127_308;
   wire [12:0] v3_1615207127_309;
   wire [12:0] v3_1615207127_310;
   wire [12:0] v3_1615207127_311;
   wire [12:0] v3_1615207127_312;
   wire [12:0] v3_1615207127_313;
   wire [6:0] v3_1615207127_314;
   wire [12:0] v3_1615207127_315;
   wire [12:0] v3_1615207127_316;
   wire [12:0] v3_1615207127_317;
   wire [12:0] v3_1615207127_318;
   wire [12:0] v3_1615207127_319;
   wire [12:0] v3_1615207127_320;
   wire [12:0] v3_1615207127_321;
   wire [12:0] v3_1615207127_322;
   wire [12:0] v3_1615207127_323;
   wire [12:0] v3_1615207127_324;
   wire [12:0] v3_1615207127_325;
   wire [12:0] v3_1615207127_326;
   wire [12:0] v3_1615207127_327;
   wire [12:0] v3_1615207127_328;
   wire [12:0] v3_1615207127_329;
   wire [12:0] v3_1615207127_330;
   wire [12:0] v3_1615207127_331;
   wire [12:0] v3_1615207127_332;
   wire [12:0] v3_1615207127_333;
   wire [12:0] v3_1615207127_334;
   wire [12:0] v3_1615207127_335;
   wire [12:0] v3_1615207127_336;
   wire [12:0] v3_1615207127_337;
   wire [12:0] v3_1615207127_338;
   wire [12:0] v3_1615207127_339;
   wire [12:0] v3_1615207127_340;
   wire [12:0] v3_1615207127_341;
   wire [12:0] v3_1615207127_342;
   wire [12:0] v3_1615207127_343;
   wire [12:0] v3_1615207127_344;
   wire [12:0] v3_1615207127_345;
   wire [12:0] v3_1615207127_346;
   wire [12:0] v3_1615207127_347;
   wire [12:0] v3_1615207127_348;
   wire [12:0] v3_1615207127_349;
   wire [12:0] v3_1615207127_350;
   wire [12:0] v3_1615207127_351;
   wire [12:0] v3_1615207127_352;
   wire [12:0] v3_1615207127_353;
   wire [12:0] v3_1615207127_354;
   wire [12:0] v3_1615207127_355;
   wire [12:0] v3_1615207127_356;
   wire [12:0] v3_1615207127_357;
   wire [12:0] v3_1615207127_358;
   wire [12:0] v3_1615207127_359;
   wire [12:0] v3_1615207127_360;
   wire [12:0] v3_1615207127_361;
   wire [12:0] v3_1615207127_362;
   wire [12:0] v3_1615207127_363;
   wire [12:0] v3_1615207127_364;
   wire [12:0] v3_1615207127_365;
   wire [12:0] v3_1615207127_366;
   wire [12:0] v3_1615207127_367;
   wire [12:0] v3_1615207127_368;
   wire [12:0] v3_1615207127_369;
   wire [12:0] v3_1615207127_370;
   wire [12:0] v3_1615207127_371;
   wire [12:0] v3_1615207127_372;
   wire [12:0] v3_1615207127_373;
   wire [12:0] v3_1615207127_374;
   wire [12:0] v3_1615207127_375;
   wire [12:0] v3_1615207127_376;
   wire [12:0] v3_1615207127_377;
   wire [12:0] v3_1615207127_378;
   wire [12:0] v3_1615207127_379;
   wire [12:0] v3_1615207127_380;
   wire v3_1615207127_381;
   wire [12:0] v3_1615207127_382;
   wire v3_1615207127_383;
   wire [12:0] v3_1615207127_384;
   wire v3_1615207127_385;
   wire [12:0] v3_1615207127_386;
   wire v3_1615207127_387;
   wire [12:0] v3_1615207127_388;
   wire [12:0] v3_1615207127_389;
   wire [12:0] v3_1615207127_390;
   wire [12:0] v3_1615207127_391;
   wire [12:0] v3_1615207127_392;
   wire [12:0] v3_1615207127_393;
   wire [12:0] v3_1615207127_394;
   wire [12:0] v3_1615207127_395;
   wire [12:0] v3_1615207127_396;
   wire [12:0] v3_1615207127_397;
   wire [12:0] v3_1615207127_398;
   wire [12:0] v3_1615207127_399;
   wire [12:0] v3_1615207127_400;
   wire [12:0] v3_1615207127_401;
   wire [12:0] v3_1615207127_402;
   wire [12:0] v3_1615207127_403;
   wire [12:0] v3_1615207127_404;
   wire [12:0] v3_1615207127_405;
   wire [12:0] v3_1615207127_406;
   wire [12:0] v3_1615207127_407;
   wire [12:0] v3_1615207127_408;
   wire [12:0] v3_1615207127_409;
   wire [12:0] v3_1615207127_410;
   wire [12:0] v3_1615207127_411;
   wire [12:0] v3_1615207127_412;
   wire [12:0] v3_1615207127_413;
   wire [12:0] v3_1615207127_414;
   wire [12:0] v3_1615207127_415;
   wire [12:0] v3_1615207127_416;
   wire [12:0] v3_1615207127_417;
   wire [12:0] v3_1615207127_418;
   wire [12:0] v3_1615207127_419;
   wire [12:0] v3_1615207127_420;
   wire [12:0] v3_1615207127_421;
   wire [12:0] v3_1615207127_422;
   wire [12:0] v3_1615207127_423;
   wire [12:0] v3_1615207127_424;
   wire [12:0] v3_1615207127_425;
   wire [12:0] v3_1615207127_426;
   wire [12:0] v3_1615207127_427;
   wire [12:0] v3_1615207127_428;
   wire [12:0] v3_1615207127_429;
   wire [12:0] v3_1615207127_430;
   wire [12:0] v3_1615207127_431;
   wire [12:0] v3_1615207127_432;
   wire [9:0] v3_1615207127_433;
   wire [12:0] v3_1615207127_434;
   wire [12:0] v3_1615207127_435;
   wire v3_1615207127_436;
   wire [12:0] v3_1615207127_437;
   wire [12:0] v3_1615207127_438;
   wire [12:0] v3_1615207127_439;
   wire [12:0] v3_1615207127_440;
   wire v3_1615207127_441;
   wire [12:0] v3_1615207127_442;
   wire [12:0] v3_1615207127_443;
   wire [12:0] v3_1615207127_444;
   wire [12:0] v3_1615207127_445;
   wire v3_1615207127_446;
   wire [12:0] v3_1615207127_447;
   wire [12:0] v3_1615207127_448;
   wire [12:0] v3_1615207127_449;
   wire [12:0] v3_1615207127_450;
   wire v3_1615207127_451;
   wire [12:0] v3_1615207127_452;
   wire [12:0] v3_1615207127_453;
   wire [5:0] v3_1615207127_454;
   wire [5:0] v3_1615207127_455;
   wire [5:0] v3_1615207127_456;
   wire [5:0] v3_1615207127_457;
   wire [5:0] v3_1615207127_458;
   wire [5:0] v3_1615207127_459;
   wire [5:0] v3_1615207127_460;
   wire [5:0] v3_1615207127_461;
   wire [5:0] v3_1615207127_462;
   wire [5:0] v3_1615207127_463;
   wire [5:0] v3_1615207127_464;
   wire [5:0] v3_1615207127_465;
   wire [5:0] v3_1615207127_466;
   wire [5:0] v3_1615207127_467;
   wire [5:0] v3_1615207127_468;
   wire [5:0] v3_1615207127_469;
   wire [5:0] v3_1615207127_470;
   wire [5:0] v3_1615207127_471;
   wire [5:0] v3_1615207127_472;
   wire [5:0] v3_1615207127_473;
   wire [5:0] v3_1615207127_474;
   wire [5:0] v3_1615207127_475;
   wire [5:0] v3_1615207127_476;
   wire [5:0] v3_1615207127_477;
   wire [5:0] v3_1615207127_478;
   wire [5:0] v3_1615207127_479;
   wire [5:0] v3_1615207127_480;
   wire [5:0] v3_1615207127_481;
   wire [5:0] v3_1615207127_482;
   wire [5:0] v3_1615207127_483;
   wire [5:0] v3_1615207127_484;
   wire v3_1615207127_485;
   wire [6:0] v3_1615207127_486;
   wire [6:0] v3_1615207127_487;
   wire [6:0] v3_1615207127_488;
   wire [6:0] v3_1615207127_489;
   wire [6:0] v3_1615207127_490;
   wire [6:0] v3_1615207127_491;
   wire [6:0] v3_1615207127_492;
   wire [5:0] v3_1615207127_493;
   wire [5:0] v3_1615207127_494;
   wire [5:0] v3_1615207127_495;
   wire [5:0] v3_1615207127_496;
   wire [5:0] v3_1615207127_497;
   wire [5:0] v3_1615207127_498;
   wire [5:0] v3_1615207127_499;
   wire [5:0] v3_1615207127_500;
   wire [5:0] v3_1615207127_501;
   wire [5:0] v3_1615207127_502;
   wire [5:0] v3_1615207127_503;
   wire [5:0] v3_1615207127_504;
   wire [5:0] v3_1615207127_505;
   wire [5:0] v3_1615207127_506;
   wire [5:0] v3_1615207127_507;
   wire [5:0] v3_1615207127_508;
   wire [5:0] v3_1615207127_509;
   wire [5:0] v3_1615207127_510;
   wire [5:0] v3_1615207127_511;
   wire [5:0] v3_1615207127_512;
   wire [5:0] v3_1615207127_513;
   wire [5:0] v3_1615207127_514;
   wire [5:0] v3_1615207127_515;
   wire [5:0] v3_1615207127_516;
   wire [5:0] v3_1615207127_517;
   wire [5:0] v3_1615207127_518;
   wire [5:0] v3_1615207127_519;
   wire [5:0] v3_1615207127_520;
   wire [5:0] v3_1615207127_521;
   wire [5:0] v3_1615207127_522;
   wire [5:0] v3_1615207127_523;
   wire [5:0] v3_1615207127_524;
   wire [5:0] v3_1615207127_525;
   wire v3_1615207127_526;
   wire [6:0] v3_1615207127_527;
   wire [6:0] v3_1615207127_528;
   wire [6:0] v3_1615207127_529;
   wire [6:0] v3_1615207127_530;
   wire [6:0] v3_1615207127_531;
   wire [6:0] v3_1615207127_532;
   wire [5:0] v3_1615207127_533;
   wire [5:0] v3_1615207127_534;
   wire [5:0] v3_1615207127_535;
   wire [5:0] v3_1615207127_536;
   wire [5:0] v3_1615207127_537;
   wire [5:0] v3_1615207127_538;
   wire [5:0] v3_1615207127_539;
   wire [5:0] v3_1615207127_540;
   wire [5:0] v3_1615207127_541;
   wire [5:0] v3_1615207127_542;
   wire [5:0] v3_1615207127_543;
   wire [5:0] v3_1615207127_544;
   wire [5:0] v3_1615207127_545;
   wire [5:0] v3_1615207127_546;
   wire [5:0] v3_1615207127_547;
   wire [5:0] v3_1615207127_548;
   wire [5:0] v3_1615207127_549;
   wire [5:0] v3_1615207127_550;
   wire [5:0] v3_1615207127_551;
   wire [5:0] v3_1615207127_552;
   wire [5:0] v3_1615207127_553;
   wire [5:0] v3_1615207127_554;
   wire [5:0] v3_1615207127_555;
   wire [5:0] v3_1615207127_556;
   wire [5:0] v3_1615207127_557;
   wire [5:0] v3_1615207127_558;
   wire [5:0] v3_1615207127_559;
   wire [5:0] v3_1615207127_560;
   wire [5:0] v3_1615207127_561;
   wire v3_1615207127_562;
   wire [6:0] v3_1615207127_563;
   wire [6:0] v3_1615207127_564;
   wire [6:0] v3_1615207127_565;
   wire [6:0] v3_1615207127_566;
   wire [6:0] v3_1615207127_567;
   wire [6:0] v3_1615207127_568;
   wire [5:0] v3_1615207127_569;
   wire [5:0] v3_1615207127_570;
   wire [5:0] v3_1615207127_571;
   wire [5:0] v3_1615207127_572;
   wire [5:0] v3_1615207127_573;
   wire [5:0] v3_1615207127_574;
   wire [5:0] v3_1615207127_575;
   wire [5:0] v3_1615207127_576;
   wire [5:0] v3_1615207127_577;
   wire [5:0] v3_1615207127_578;
   wire [5:0] v3_1615207127_579;
   wire [5:0] v3_1615207127_580;
   wire [5:0] v3_1615207127_581;
   wire [5:0] v3_1615207127_582;
   wire [5:0] v3_1615207127_583;
   wire [5:0] v3_1615207127_584;
   wire [5:0] v3_1615207127_585;
   wire [5:0] v3_1615207127_586;
   wire [5:0] v3_1615207127_587;
   wire [5:0] v3_1615207127_588;
   wire [5:0] v3_1615207127_589;
   wire [5:0] v3_1615207127_590;
   wire [5:0] v3_1615207127_591;
   wire [5:0] v3_1615207127_592;
   wire [5:0] v3_1615207127_593;
   wire [5:0] v3_1615207127_594;
   wire [5:0] v3_1615207127_595;
   wire [5:0] v3_1615207127_596;
   wire [5:0] v3_1615207127_597;
   wire [5:0] v3_1615207127_598;
   wire [5:0] v3_1615207127_599;
   wire [5:0] v3_1615207127_600;
   wire [5:0] v3_1615207127_601;
   wire v3_1615207127_602;
   wire [6:0] v3_1615207127_603;
   wire [6:0] v3_1615207127_604;
   wire [6:0] v3_1615207127_605;
   wire [6:0] v3_1615207127_606;
   wire [6:0] v3_1615207127_607;
   wire [6:0] v3_1615207127_608;
   wire [5:0] v3_1615207127_609;
   wire [5:0] v3_1615207127_610;
   wire [5:0] v3_1615207127_611;

   // Output Net Declarations
   wire [5:0] coinOutA;
   wire [5:0] coinOutB;
   wire [5:0] coinOutC;
   wire [5:0] coinOutD;
   wire [1:0] itemTypeOut;
   wire [2:0] itemNumberOut;
   wire [1:0] serviceTypeOut;

   // Combinational Assignments
   assign v3_1615207127_0 = 1'b0; 
   assign v3_1615207127_27 = v3_1615207127_75 ? v3_1615207127_74 : v3_1615207127_28;
   assign v3_1615207127_28 = v3_1615207127_17 ? v3_1615207127_30 : v3_1615207127_29;
   assign v3_1615207127_29 = v3_1615207127_10;
   assign v3_1615207127_30 = v3_1615207127_73 ? v3_1615207127_67 : v3_1615207127_31;
   assign v3_1615207127_31 = v3_1615207127_66 ? v3_1615207127_65 : v3_1615207127_32;
   assign v3_1615207127_32 = v3_1615207127_64 ? v3_1615207127_63 : v3_1615207127_33;
   assign v3_1615207127_33 = v3_1615207127_61 ? v3_1615207127_51 : v3_1615207127_34;
   assign v3_1615207127_34 = v3_1615207127_49 ? v3_1615207127_48 : v3_1615207127_35;
   assign v3_1615207127_35 = v3_1615207127_46 ? v3_1615207127_45 : v3_1615207127_36;
   assign v3_1615207127_36 = v3_1615207127_43 ? v3_1615207127_38 : v3_1615207127_37;
   assign v3_1615207127_37 = v3_1615207127_10;
   assign v3_1615207127_38 = v3_1615207127_42 ? v3_1615207127_40 : v3_1615207127_39;
   assign v3_1615207127_39 = v3_1615207127_10;
   assign v3_1615207127_40 = v3_1615207127_41;
   assign v3_1615207127_41 = 6'b000000; 
   assign v3_1615207127_42 = v3_1615207127_25 == v3_1615207127_41;
   assign v3_1615207127_43 = v3_1615207127_22 >= v3_1615207127_44;
   assign v3_1615207127_44 = 13'b00000_00000001; 
   assign v3_1615207127_45 = v3_1615207127_10;
   assign v3_1615207127_46 = v3_1615207127_19 == v3_1615207127_47;
   assign v3_1615207127_47 = 2'b10; 
   assign v3_1615207127_48 = v3_1615207127_10;
   assign v3_1615207127_49 = v3_1615207127_19 == v3_1615207127_50;
   assign v3_1615207127_50 = 2'b01; 
   assign v3_1615207127_51 = v3_1615207127_59 ? v3_1615207127_53 : v3_1615207127_52;
   assign v3_1615207127_52 = v3_1615207127_10;
   assign v3_1615207127_53 = v3_1615207127_58 ? v3_1615207127_57 : v3_1615207127_54;
   assign v3_1615207127_54 = v3_1615207127_56;
   assign v3_1615207127_55 = 6'b000001; 
   assign v3_1615207127_56 = v3_1615207127_10 + v3_1615207127_55;
   assign v3_1615207127_57 = v3_1615207127_10;
   assign v3_1615207127_58 = v3_1615207127_23 == v3_1615207127_41;
   assign v3_1615207127_59 = v3_1615207127_22 >= v3_1615207127_60;
   assign v3_1615207127_60 = 13'b00000_00110010; 
   assign v3_1615207127_61 = v3_1615207127_19 == v3_1615207127_62;
   assign v3_1615207127_62 = 2'b00; 
   assign v3_1615207127_63 = v3_1615207127_10;
   assign v3_1615207127_64 = ~v3_1615207127_18;
   assign v3_1615207127_65 = v3_1615207127_10;
   assign v3_1615207127_66 = v3_1615207127_16 == v3_1615207127_62;
   assign v3_1615207127_67 = v3_1615207127_70 ? v3_1615207127_69 : v3_1615207127_68;
   assign v3_1615207127_68 = v3_1615207127_10;
   assign v3_1615207127_69 = v3_1615207127_41;
   assign v3_1615207127_70 = ~v3_1615207127_71;
   assign v3_1615207127_71 = itemNumberIn == v3_1615207127_72;
   assign v3_1615207127_72 = 3'b000; 
   assign v3_1615207127_73 = v3_1615207127_16 == v3_1615207127_50;
   assign v3_1615207127_74 = v3_1615207127_41;
   assign v3_1615207127_75 = ~reset;
   assign v3_1615207127_76 = 6'b000000; 
   assign v3_1615207127_77 = v3_1615207127_75 ? v3_1615207127_107 : v3_1615207127_78;
   assign v3_1615207127_78 = v3_1615207127_17 ? v3_1615207127_80 : v3_1615207127_79;
   assign v3_1615207127_79 = v3_1615207127_11;
   assign v3_1615207127_80 = v3_1615207127_73 ? v3_1615207127_104 : v3_1615207127_81;
   assign v3_1615207127_81 = v3_1615207127_66 ? v3_1615207127_103 : v3_1615207127_82;
   assign v3_1615207127_82 = v3_1615207127_64 ? v3_1615207127_102 : v3_1615207127_83;
   assign v3_1615207127_83 = v3_1615207127_61 ? v3_1615207127_101 : v3_1615207127_84;
   assign v3_1615207127_84 = v3_1615207127_49 ? v3_1615207127_92 : v3_1615207127_85;
   assign v3_1615207127_85 = v3_1615207127_46 ? v3_1615207127_91 : v3_1615207127_86;
   assign v3_1615207127_86 = v3_1615207127_43 ? v3_1615207127_88 : v3_1615207127_87;
   assign v3_1615207127_87 = v3_1615207127_11;
   assign v3_1615207127_88 = v3_1615207127_42 ? v3_1615207127_90 : v3_1615207127_89;
   assign v3_1615207127_89 = v3_1615207127_11;
   assign v3_1615207127_90 = v3_1615207127_41;
   assign v3_1615207127_91 = v3_1615207127_11;
   assign v3_1615207127_92 = v3_1615207127_99 ? v3_1615207127_94 : v3_1615207127_93;
   assign v3_1615207127_93 = v3_1615207127_11;
   assign v3_1615207127_94 = v3_1615207127_98 ? v3_1615207127_97 : v3_1615207127_95;
   assign v3_1615207127_95 = v3_1615207127_96;
   assign v3_1615207127_96 = v3_1615207127_11 + v3_1615207127_55;
   assign v3_1615207127_97 = v3_1615207127_11;
   assign v3_1615207127_98 = v3_1615207127_24 == v3_1615207127_41;
   assign v3_1615207127_99 = v3_1615207127_22 >= v3_1615207127_100;
   assign v3_1615207127_100 = 13'b00000_00001010; 
   assign v3_1615207127_101 = v3_1615207127_11;
   assign v3_1615207127_102 = v3_1615207127_11;
   assign v3_1615207127_103 = v3_1615207127_11;
   assign v3_1615207127_104 = v3_1615207127_70 ? v3_1615207127_106 : v3_1615207127_105;
   assign v3_1615207127_105 = v3_1615207127_11;
   assign v3_1615207127_106 = v3_1615207127_41;
   assign v3_1615207127_107 = v3_1615207127_41;
   assign v3_1615207127_108 = 6'b000000; 
   assign v3_1615207127_109 = v3_1615207127_75 ? v3_1615207127_139 : v3_1615207127_110;
   assign v3_1615207127_110 = v3_1615207127_17 ? v3_1615207127_112 : v3_1615207127_111;
   assign v3_1615207127_111 = v3_1615207127_12;
   assign v3_1615207127_112 = v3_1615207127_73 ? v3_1615207127_136 : v3_1615207127_113;
   assign v3_1615207127_113 = v3_1615207127_66 ? v3_1615207127_135 : v3_1615207127_114;
   assign v3_1615207127_114 = v3_1615207127_64 ? v3_1615207127_134 : v3_1615207127_115;
   assign v3_1615207127_115 = v3_1615207127_61 ? v3_1615207127_133 : v3_1615207127_116;
   assign v3_1615207127_116 = v3_1615207127_49 ? v3_1615207127_132 : v3_1615207127_117;
   assign v3_1615207127_117 = v3_1615207127_46 ? v3_1615207127_123 : v3_1615207127_118;
   assign v3_1615207127_118 = v3_1615207127_43 ? v3_1615207127_120 : v3_1615207127_119;
   assign v3_1615207127_119 = v3_1615207127_12;
   assign v3_1615207127_120 = v3_1615207127_42 ? v3_1615207127_122 : v3_1615207127_121;
   assign v3_1615207127_121 = v3_1615207127_12;
   assign v3_1615207127_122 = v3_1615207127_41;
   assign v3_1615207127_123 = v3_1615207127_130 ? v3_1615207127_125 : v3_1615207127_124;
   assign v3_1615207127_124 = v3_1615207127_12;
   assign v3_1615207127_125 = v3_1615207127_129 ? v3_1615207127_128 : v3_1615207127_126;
   assign v3_1615207127_126 = v3_1615207127_127;
   assign v3_1615207127_127 = v3_1615207127_12 + v3_1615207127_55;
   assign v3_1615207127_128 = v3_1615207127_12;
   assign v3_1615207127_129 = v3_1615207127_26 == v3_1615207127_41;
   assign v3_1615207127_130 = v3_1615207127_22 >= v3_1615207127_131;
   assign v3_1615207127_131 = 13'b00000_00000101; 
   assign v3_1615207127_132 = v3_1615207127_12;
   assign v3_1615207127_133 = v3_1615207127_12;
   assign v3_1615207127_134 = v3_1615207127_12;
   assign v3_1615207127_135 = v3_1615207127_12;
   assign v3_1615207127_136 = v3_1615207127_70 ? v3_1615207127_138 : v3_1615207127_137;
   assign v3_1615207127_137 = v3_1615207127_12;
   assign v3_1615207127_138 = v3_1615207127_41;
   assign v3_1615207127_139 = v3_1615207127_41;
   assign v3_1615207127_140 = 6'b000000; 
   assign v3_1615207127_141 = v3_1615207127_75 ? v3_1615207127_164 : v3_1615207127_142;
   assign v3_1615207127_142 = v3_1615207127_17 ? v3_1615207127_144 : v3_1615207127_143;
   assign v3_1615207127_143 = v3_1615207127_13;
   assign v3_1615207127_144 = v3_1615207127_73 ? v3_1615207127_161 : v3_1615207127_145;
   assign v3_1615207127_145 = v3_1615207127_66 ? v3_1615207127_160 : v3_1615207127_146;
   assign v3_1615207127_146 = v3_1615207127_64 ? v3_1615207127_159 : v3_1615207127_147;
   assign v3_1615207127_147 = v3_1615207127_61 ? v3_1615207127_158 : v3_1615207127_148;
   assign v3_1615207127_148 = v3_1615207127_49 ? v3_1615207127_157 : v3_1615207127_149;
   assign v3_1615207127_149 = v3_1615207127_46 ? v3_1615207127_156 : v3_1615207127_150;
   assign v3_1615207127_150 = v3_1615207127_43 ? v3_1615207127_152 : v3_1615207127_151;
   assign v3_1615207127_151 = v3_1615207127_13;
   assign v3_1615207127_152 = v3_1615207127_42 ? v3_1615207127_155 : v3_1615207127_153;
   assign v3_1615207127_153 = v3_1615207127_154;
   assign v3_1615207127_154 = v3_1615207127_13 + v3_1615207127_55;
   assign v3_1615207127_155 = v3_1615207127_41;
   assign v3_1615207127_156 = v3_1615207127_13;
   assign v3_1615207127_157 = v3_1615207127_13;
   assign v3_1615207127_158 = v3_1615207127_13;
   assign v3_1615207127_159 = v3_1615207127_13;
   assign v3_1615207127_160 = v3_1615207127_13;
   assign v3_1615207127_161 = v3_1615207127_70 ? v3_1615207127_163 : v3_1615207127_162;
   assign v3_1615207127_162 = v3_1615207127_13;
   assign v3_1615207127_163 = v3_1615207127_41;
   assign v3_1615207127_164 = v3_1615207127_41;
   assign v3_1615207127_165 = 6'b000000; 
   assign v3_1615207127_166 = v3_1615207127_75 ? v3_1615207127_174 : v3_1615207127_167;
   assign v3_1615207127_167 = v3_1615207127_17 ? v3_1615207127_169 : v3_1615207127_168;
   assign v3_1615207127_168 = v3_1615207127_14;
   assign v3_1615207127_169 = v3_1615207127_73 ? v3_1615207127_171 : v3_1615207127_170;
   assign v3_1615207127_170 = v3_1615207127_14;
   assign v3_1615207127_171 = v3_1615207127_70 ? v3_1615207127_173 : v3_1615207127_172;
   assign v3_1615207127_172 = v3_1615207127_14;
   assign v3_1615207127_173 = itemTypeIn;
   assign v3_1615207127_174 = v3_1615207127_62;
   assign v3_1615207127_175 = 2'b00; 
   assign v3_1615207127_176 = v3_1615207127_75 ? v3_1615207127_207 : v3_1615207127_177;
   assign v3_1615207127_177 = v3_1615207127_17 ? v3_1615207127_179 : v3_1615207127_178;
   assign v3_1615207127_178 = v3_1615207127_15;
   assign v3_1615207127_179 = v3_1615207127_73 ? v3_1615207127_204 : v3_1615207127_180;
   assign v3_1615207127_180 = v3_1615207127_66 ? v3_1615207127_203 : v3_1615207127_181;
   assign v3_1615207127_181 = v3_1615207127_64 ? v3_1615207127_197 : v3_1615207127_182;
   assign v3_1615207127_182 = v3_1615207127_61 ? v3_1615207127_196 : v3_1615207127_183;
   assign v3_1615207127_183 = v3_1615207127_49 ? v3_1615207127_195 : v3_1615207127_184;
   assign v3_1615207127_184 = v3_1615207127_46 ? v3_1615207127_194 : v3_1615207127_185;
   assign v3_1615207127_185 = v3_1615207127_43 ? v3_1615207127_187 : v3_1615207127_186;
   assign v3_1615207127_186 = v3_1615207127_15;
   assign v3_1615207127_187 = v3_1615207127_42 ? v3_1615207127_189 : v3_1615207127_188;
   assign v3_1615207127_188 = v3_1615207127_15;
   assign v3_1615207127_189 = v3_1615207127_20 ? v3_1615207127_191 : v3_1615207127_190;
   assign v3_1615207127_190 = v3_1615207127_72;
   assign v3_1615207127_191 = v3_1615207127_193;
   assign v3_1615207127_192 = 3'b001; 
   assign v3_1615207127_193 = v3_1615207127_15 - v3_1615207127_192;
   assign v3_1615207127_194 = v3_1615207127_15;
   assign v3_1615207127_195 = v3_1615207127_15;
   assign v3_1615207127_196 = v3_1615207127_15;
   assign v3_1615207127_197 = v3_1615207127_201 ? v3_1615207127_199 : v3_1615207127_198;
   assign v3_1615207127_198 = v3_1615207127_15;
   assign v3_1615207127_199 = v3_1615207127_20 ? v3_1615207127_191 : v3_1615207127_200;
   assign v3_1615207127_200 = v3_1615207127_72;
   assign v3_1615207127_201 = ~v3_1615207127_202;
   assign v3_1615207127_202 = v3_1615207127_21 >= v3_1615207127_22;
   assign v3_1615207127_203 = v3_1615207127_15;
   assign v3_1615207127_204 = v3_1615207127_70 ? v3_1615207127_206 : v3_1615207127_205;
   assign v3_1615207127_205 = v3_1615207127_15;
   assign v3_1615207127_206 = itemNumberIn;
   assign v3_1615207127_207 = v3_1615207127_72;
   assign v3_1615207127_208 = 3'b000; 
   assign v3_1615207127_209 = v3_1615207127_75 ? v3_1615207127_229 : v3_1615207127_210;
   assign v3_1615207127_210 = v3_1615207127_17 ? v3_1615207127_212 : v3_1615207127_211;
   assign v3_1615207127_211 = v3_1615207127_16;
   assign v3_1615207127_212 = v3_1615207127_73 ? v3_1615207127_226 : v3_1615207127_213;
   assign v3_1615207127_213 = v3_1615207127_66 ? v3_1615207127_225 : v3_1615207127_214;
   assign v3_1615207127_214 = v3_1615207127_64 ? v3_1615207127_224 : v3_1615207127_215;
   assign v3_1615207127_215 = v3_1615207127_61 ? v3_1615207127_223 : v3_1615207127_216;
   assign v3_1615207127_216 = v3_1615207127_49 ? v3_1615207127_222 : v3_1615207127_217;
   assign v3_1615207127_217 = v3_1615207127_46 ? v3_1615207127_221 : v3_1615207127_218;
   assign v3_1615207127_218 = v3_1615207127_43 ? v3_1615207127_220 : v3_1615207127_219;
   assign v3_1615207127_219 = v3_1615207127_62;
   assign v3_1615207127_220 = v3_1615207127_16;
   assign v3_1615207127_221 = v3_1615207127_16;
   assign v3_1615207127_222 = v3_1615207127_16;
   assign v3_1615207127_223 = v3_1615207127_16;
   assign v3_1615207127_224 = v3_1615207127_16;
   assign v3_1615207127_225 = v3_1615207127_50;
   assign v3_1615207127_226 = v3_1615207127_70 ? v3_1615207127_228 : v3_1615207127_227;
   assign v3_1615207127_227 = v3_1615207127_16;
   assign v3_1615207127_228 = v3_1615207127_47;
   assign v3_1615207127_229 = v3_1615207127_50;
   assign v3_1615207127_230 = 2'b00; 
   assign v3_1615207127_231 = v3_1615207127_75 ? v3_1615207127_233 : v3_1615207127_232;
   assign v3_1615207127_232 = v3_1615207127_17;
   assign v3_1615207127_233 = v3_1615207127_234;
   assign v3_1615207127_234 = 1'b1; 
   assign v3_1615207127_235 = 1'b0; 
   assign v3_1615207127_236 = v3_1615207127_75 ? v3_1615207127_253 : v3_1615207127_237;
   assign v3_1615207127_237 = v3_1615207127_17 ? v3_1615207127_239 : v3_1615207127_238;
   assign v3_1615207127_238 = v3_1615207127_18;
   assign v3_1615207127_239 = v3_1615207127_73 ? v3_1615207127_249 : v3_1615207127_240;
   assign v3_1615207127_240 = v3_1615207127_66 ? v3_1615207127_248 : v3_1615207127_241;
   assign v3_1615207127_241 = v3_1615207127_64 ? v3_1615207127_243 : v3_1615207127_242;
   assign v3_1615207127_242 = v3_1615207127_18;
   assign v3_1615207127_243 = v3_1615207127_201 ? v3_1615207127_245 : v3_1615207127_244;
   assign v3_1615207127_244 = v3_1615207127_234;
   assign v3_1615207127_245 = v3_1615207127_20 ? v3_1615207127_247 : v3_1615207127_246;
   assign v3_1615207127_246 = v3_1615207127_234;
   assign v3_1615207127_247 = v3_1615207127_18;
   assign v3_1615207127_248 = v3_1615207127_18;
   assign v3_1615207127_249 = v3_1615207127_70 ? v3_1615207127_251 : v3_1615207127_250;
   assign v3_1615207127_250 = v3_1615207127_18;
   assign v3_1615207127_251 = v3_1615207127_252;
   assign v3_1615207127_252 = 1'b0; 
   assign v3_1615207127_253 = v3_1615207127_252;
   assign v3_1615207127_254 = 1'b0; 
   assign v3_1615207127_255 = v3_1615207127_75 ? v3_1615207127_290 : v3_1615207127_256;
   assign v3_1615207127_256 = v3_1615207127_17 ? v3_1615207127_258 : v3_1615207127_257;
   assign v3_1615207127_257 = v3_1615207127_19;
   assign v3_1615207127_258 = v3_1615207127_73 ? v3_1615207127_287 : v3_1615207127_259;
   assign v3_1615207127_259 = v3_1615207127_66 ? v3_1615207127_286 : v3_1615207127_260;
   assign v3_1615207127_260 = v3_1615207127_64 ? v3_1615207127_285 : v3_1615207127_261;
   assign v3_1615207127_261 = v3_1615207127_61 ? v3_1615207127_280 : v3_1615207127_262;
   assign v3_1615207127_262 = v3_1615207127_49 ? v3_1615207127_275 : v3_1615207127_263;
   assign v3_1615207127_263 = v3_1615207127_46 ? v3_1615207127_269 : v3_1615207127_264;
   assign v3_1615207127_264 = v3_1615207127_43 ? v3_1615207127_266 : v3_1615207127_265;
   assign v3_1615207127_265 = v3_1615207127_19;
   assign v3_1615207127_266 = v3_1615207127_42 ? v3_1615207127_268 : v3_1615207127_267;
   assign v3_1615207127_267 = v3_1615207127_19;
   assign v3_1615207127_268 = v3_1615207127_62;
   assign v3_1615207127_269 = v3_1615207127_130 ? v3_1615207127_272 : v3_1615207127_270;
   assign v3_1615207127_270 = v3_1615207127_271;
   assign v3_1615207127_271 = 2'b11; 
   assign v3_1615207127_272 = v3_1615207127_129 ? v3_1615207127_274 : v3_1615207127_273;
   assign v3_1615207127_273 = v3_1615207127_19;
   assign v3_1615207127_274 = v3_1615207127_271;
   assign v3_1615207127_275 = v3_1615207127_99 ? v3_1615207127_277 : v3_1615207127_276;
   assign v3_1615207127_276 = v3_1615207127_47;
   assign v3_1615207127_277 = v3_1615207127_98 ? v3_1615207127_279 : v3_1615207127_278;
   assign v3_1615207127_278 = v3_1615207127_19;
   assign v3_1615207127_279 = v3_1615207127_47;
   assign v3_1615207127_280 = v3_1615207127_59 ? v3_1615207127_282 : v3_1615207127_281;
   assign v3_1615207127_281 = v3_1615207127_50;
   assign v3_1615207127_282 = v3_1615207127_58 ? v3_1615207127_284 : v3_1615207127_283;
   assign v3_1615207127_283 = v3_1615207127_19;
   assign v3_1615207127_284 = v3_1615207127_50;
   assign v3_1615207127_285 = v3_1615207127_19;
   assign v3_1615207127_286 = v3_1615207127_19;
   assign v3_1615207127_287 = v3_1615207127_70 ? v3_1615207127_289 : v3_1615207127_288;
   assign v3_1615207127_288 = v3_1615207127_19;
   assign v3_1615207127_289 = v3_1615207127_62;
   assign v3_1615207127_290 = v3_1615207127_62;
   assign v3_1615207127_291 = 2'b00; 
   assign v3_1615207127_292 = v3_1615207127_75 ? v3_1615207127_300 : v3_1615207127_293;
   assign v3_1615207127_293 = v3_1615207127_17 ? v3_1615207127_295 : v3_1615207127_294;
   assign v3_1615207127_294 = v3_1615207127_20;
   assign v3_1615207127_295 = v3_1615207127_73 ? v3_1615207127_297 : v3_1615207127_296;
   assign v3_1615207127_296 = v3_1615207127_20;
   assign v3_1615207127_297 = v3_1615207127_70 ? v3_1615207127_299 : v3_1615207127_298;
   assign v3_1615207127_298 = v3_1615207127_20;
   assign v3_1615207127_299 = forceIn;
   assign v3_1615207127_300 = v3_1615207127_252;
   assign v3_1615207127_301 = 1'b0; 
   assign v3_1615207127_302 = v3_1615207127_75 ? v3_1615207127_332 : v3_1615207127_303;
   assign v3_1615207127_303 = v3_1615207127_17 ? v3_1615207127_305 : v3_1615207127_304;
   assign v3_1615207127_304 = v3_1615207127_21;
   assign v3_1615207127_305 = v3_1615207127_73 ? v3_1615207127_307 : v3_1615207127_306;
   assign v3_1615207127_306 = v3_1615207127_21;
   assign v3_1615207127_307 = v3_1615207127_70 ? v3_1615207127_309 : v3_1615207127_308;
   assign v3_1615207127_308 = v3_1615207127_21;
   assign v3_1615207127_309 = v3_1615207127_331;
   assign v3_1615207127_310 = v3_1615207127_326;
   assign v3_1615207127_311 = v3_1615207127_321;
   assign v3_1615207127_312 = v3_1615207127_316;
   assign v3_1615207127_313 = v3_1615207127_315;
   assign v3_1615207127_314 = 7'b0000000; 
   assign v3_1615207127_315 = {v3_1615207127_314, coinInA};
   assign v3_1615207127_316 = v3_1615207127_60 * v3_1615207127_313;
   assign v3_1615207127_317 = v3_1615207127_320;
   assign v3_1615207127_318 = v3_1615207127_319;
   assign v3_1615207127_319 = {v3_1615207127_314, coinInB};
   assign v3_1615207127_320 = v3_1615207127_100 * v3_1615207127_318;
   assign v3_1615207127_321 = v3_1615207127_312 + v3_1615207127_317;
   assign v3_1615207127_322 = v3_1615207127_325;
   assign v3_1615207127_323 = v3_1615207127_324;
   assign v3_1615207127_324 = {v3_1615207127_314, coinInC};
   assign v3_1615207127_325 = v3_1615207127_131 * v3_1615207127_323;
   assign v3_1615207127_326 = v3_1615207127_311 + v3_1615207127_322;
   assign v3_1615207127_327 = v3_1615207127_330;
   assign v3_1615207127_328 = v3_1615207127_329;
   assign v3_1615207127_329 = {v3_1615207127_314, coinInD};
   assign v3_1615207127_330 = v3_1615207127_44 * v3_1615207127_328;
   assign v3_1615207127_331 = v3_1615207127_310 + v3_1615207127_327;
   assign v3_1615207127_332 = v3_1615207127_333;
   assign v3_1615207127_333 = 13'b00000_00000000; 
   assign v3_1615207127_334 = 13'b00000_00000000; 
   assign v3_1615207127_335 = v3_1615207127_75 ? v3_1615207127_452 : v3_1615207127_336;
   assign v3_1615207127_336 = v3_1615207127_17 ? v3_1615207127_338 : v3_1615207127_337;
   assign v3_1615207127_337 = v3_1615207127_22;
   assign v3_1615207127_338 = v3_1615207127_73 ? v3_1615207127_425 : v3_1615207127_339;
   assign v3_1615207127_339 = v3_1615207127_66 ? v3_1615207127_424 : v3_1615207127_340;
   assign v3_1615207127_340 = v3_1615207127_64 ? v3_1615207127_407 : v3_1615207127_341;
   assign v3_1615207127_341 = v3_1615207127_61 ? v3_1615207127_401 : v3_1615207127_342;
   assign v3_1615207127_342 = v3_1615207127_49 ? v3_1615207127_395 : v3_1615207127_343;
   assign v3_1615207127_343 = v3_1615207127_46 ? v3_1615207127_389 : v3_1615207127_344;
   assign v3_1615207127_344 = v3_1615207127_43 ? v3_1615207127_346 : v3_1615207127_345;
   assign v3_1615207127_345 = v3_1615207127_22;
   assign v3_1615207127_346 = v3_1615207127_42 ? v3_1615207127_349 : v3_1615207127_347;
   assign v3_1615207127_347 = v3_1615207127_348;
   assign v3_1615207127_348 = v3_1615207127_22 - v3_1615207127_44;
   assign v3_1615207127_349 = v3_1615207127_20 ? v3_1615207127_351 : v3_1615207127_350;
   assign v3_1615207127_350 = v3_1615207127_21;
   assign v3_1615207127_351 = v3_1615207127_388;
   assign v3_1615207127_352 = v3_1615207127_375;
   assign v3_1615207127_353 = v3_1615207127_374;
   assign v3_1615207127_354 = v3_1615207127_369;
   assign v3_1615207127_355 = v3_1615207127_364;
   assign v3_1615207127_356 = v3_1615207127_359;
   assign v3_1615207127_357 = v3_1615207127_358;
   assign v3_1615207127_358 = {v3_1615207127_314, v3_1615207127_10};
   assign v3_1615207127_359 = v3_1615207127_60 * v3_1615207127_357;
   assign v3_1615207127_360 = v3_1615207127_363;
   assign v3_1615207127_361 = v3_1615207127_362;
   assign v3_1615207127_362 = {v3_1615207127_314, v3_1615207127_11};
   assign v3_1615207127_363 = v3_1615207127_100 * v3_1615207127_361;
   assign v3_1615207127_364 = v3_1615207127_356 + v3_1615207127_360;
   assign v3_1615207127_365 = v3_1615207127_368;
   assign v3_1615207127_366 = v3_1615207127_367;
   assign v3_1615207127_367 = {v3_1615207127_314, v3_1615207127_12};
   assign v3_1615207127_368 = v3_1615207127_131 * v3_1615207127_366;
   assign v3_1615207127_369 = v3_1615207127_355 + v3_1615207127_365;
   assign v3_1615207127_370 = v3_1615207127_373;
   assign v3_1615207127_371 = v3_1615207127_372;
   assign v3_1615207127_372 = {v3_1615207127_314, v3_1615207127_13};
   assign v3_1615207127_373 = v3_1615207127_44 * v3_1615207127_371;
   assign v3_1615207127_374 = v3_1615207127_354 + v3_1615207127_370;
   assign v3_1615207127_375 = v3_1615207127_353 + v3_1615207127_22;
   assign v3_1615207127_376 = v3_1615207127_387 ? v3_1615207127_386 : v3_1615207127_377;
   assign v3_1615207127_377 = v3_1615207127_385 ? v3_1615207127_384 : v3_1615207127_378;
   assign v3_1615207127_378 = v3_1615207127_383 ? v3_1615207127_382 : v3_1615207127_379;
   assign v3_1615207127_379 = v3_1615207127_381 ? v3_1615207127_380 : v3_1615207127_333;
   assign v3_1615207127_380 = 13'b00000_01100100; 
   assign v3_1615207127_381 = v3_1615207127_14 == v3_1615207127_271;
   assign v3_1615207127_382 = 13'b00000_01001011; 
   assign v3_1615207127_383 = v3_1615207127_14 == v3_1615207127_47;
   assign v3_1615207127_384 = 13'b00000_00011001; 
   assign v3_1615207127_385 = v3_1615207127_14 == v3_1615207127_50;
   assign v3_1615207127_386 = 13'b00000_00001111; 
   assign v3_1615207127_387 = v3_1615207127_14 == v3_1615207127_62;
   assign v3_1615207127_388 = v3_1615207127_352 + v3_1615207127_376;
   assign v3_1615207127_389 = v3_1615207127_130 ? v3_1615207127_391 : v3_1615207127_390;
   assign v3_1615207127_390 = v3_1615207127_22;
   assign v3_1615207127_391 = v3_1615207127_129 ? v3_1615207127_394 : v3_1615207127_392;
   assign v3_1615207127_392 = v3_1615207127_393;
   assign v3_1615207127_393 = v3_1615207127_22 - v3_1615207127_131;
   assign v3_1615207127_394 = v3_1615207127_22;
   assign v3_1615207127_395 = v3_1615207127_99 ? v3_1615207127_397 : v3_1615207127_396;
   assign v3_1615207127_396 = v3_1615207127_22;
   assign v3_1615207127_397 = v3_1615207127_98 ? v3_1615207127_400 : v3_1615207127_398;
   assign v3_1615207127_398 = v3_1615207127_399;
   assign v3_1615207127_399 = v3_1615207127_22 - v3_1615207127_100;
   assign v3_1615207127_400 = v3_1615207127_22;
   assign v3_1615207127_401 = v3_1615207127_59 ? v3_1615207127_403 : v3_1615207127_402;
   assign v3_1615207127_402 = v3_1615207127_22;
   assign v3_1615207127_403 = v3_1615207127_58 ? v3_1615207127_406 : v3_1615207127_404;
   assign v3_1615207127_404 = v3_1615207127_405;
   assign v3_1615207127_405 = v3_1615207127_22 - v3_1615207127_60;
   assign v3_1615207127_406 = v3_1615207127_22;
   assign v3_1615207127_407 = v3_1615207127_201 ? v3_1615207127_410 : v3_1615207127_408;
   assign v3_1615207127_408 = v3_1615207127_409;
   assign v3_1615207127_409 = v3_1615207127_21 - v3_1615207127_22;
   assign v3_1615207127_410 = v3_1615207127_20 ? v3_1615207127_412 : v3_1615207127_411;
   assign v3_1615207127_411 = v3_1615207127_21;
   assign v3_1615207127_412 = v3_1615207127_387 ? v3_1615207127_422 : v3_1615207127_413;
   assign v3_1615207127_413 = v3_1615207127_385 ? v3_1615207127_420 : v3_1615207127_414;
   assign v3_1615207127_414 = v3_1615207127_383 ? v3_1615207127_418 : v3_1615207127_415;
   assign v3_1615207127_415 = v3_1615207127_381 ? v3_1615207127_416 : v3_1615207127_333;
   assign v3_1615207127_416 = v3_1615207127_417;
   assign v3_1615207127_417 = v3_1615207127_22 - v3_1615207127_380;
   assign v3_1615207127_418 = v3_1615207127_419;
   assign v3_1615207127_419 = v3_1615207127_22 - v3_1615207127_382;
   assign v3_1615207127_420 = v3_1615207127_421;
   assign v3_1615207127_421 = v3_1615207127_22 - v3_1615207127_384;
   assign v3_1615207127_422 = v3_1615207127_423;
   assign v3_1615207127_423 = v3_1615207127_22 - v3_1615207127_386;
   assign v3_1615207127_424 = v3_1615207127_22;
   assign v3_1615207127_425 = v3_1615207127_70 ? v3_1615207127_427 : v3_1615207127_426;
   assign v3_1615207127_426 = v3_1615207127_22;
   assign v3_1615207127_427 = v3_1615207127_451 ? v3_1615207127_447 : v3_1615207127_428;
   assign v3_1615207127_428 = v3_1615207127_446 ? v3_1615207127_442 : v3_1615207127_429;
   assign v3_1615207127_429 = v3_1615207127_441 ? v3_1615207127_437 : v3_1615207127_430;
   assign v3_1615207127_430 = v3_1615207127_436 ? v3_1615207127_431 : v3_1615207127_333;
   assign v3_1615207127_431 = v3_1615207127_435;
   assign v3_1615207127_432 = v3_1615207127_434;
   assign v3_1615207127_433 = 10'b00_00000000; 
   assign v3_1615207127_434 = {v3_1615207127_433, itemNumberIn};
   assign v3_1615207127_435 = v3_1615207127_432 * v3_1615207127_380;
   assign v3_1615207127_436 = itemTypeIn == v3_1615207127_271;
   assign v3_1615207127_437 = v3_1615207127_440;
   assign v3_1615207127_438 = v3_1615207127_439;
   assign v3_1615207127_439 = {v3_1615207127_433, itemNumberIn};
   assign v3_1615207127_440 = v3_1615207127_438 * v3_1615207127_382;
   assign v3_1615207127_441 = itemTypeIn == v3_1615207127_47;
   assign v3_1615207127_442 = v3_1615207127_445;
   assign v3_1615207127_443 = v3_1615207127_444;
   assign v3_1615207127_444 = {v3_1615207127_433, itemNumberIn};
   assign v3_1615207127_445 = v3_1615207127_443 * v3_1615207127_384;
   assign v3_1615207127_446 = itemTypeIn == v3_1615207127_50;
   assign v3_1615207127_447 = v3_1615207127_450;
   assign v3_1615207127_448 = v3_1615207127_449;
   assign v3_1615207127_449 = {v3_1615207127_433, itemNumberIn};
   assign v3_1615207127_450 = v3_1615207127_448 * v3_1615207127_386;
   assign v3_1615207127_451 = itemTypeIn == v3_1615207127_62;
   assign v3_1615207127_452 = v3_1615207127_333;
   assign v3_1615207127_453 = 13'b00000_00000000; 
   assign v3_1615207127_454 = v3_1615207127_75 ? v3_1615207127_493 : v3_1615207127_455;
   assign v3_1615207127_455 = v3_1615207127_17 ? v3_1615207127_457 : v3_1615207127_456;
   assign v3_1615207127_456 = v3_1615207127_23;
   assign v3_1615207127_457 = v3_1615207127_73 ? v3_1615207127_479 : v3_1615207127_458;
   assign v3_1615207127_458 = v3_1615207127_66 ? v3_1615207127_478 : v3_1615207127_459;
   assign v3_1615207127_459 = v3_1615207127_64 ? v3_1615207127_477 : v3_1615207127_460;
   assign v3_1615207127_460 = v3_1615207127_61 ? v3_1615207127_471 : v3_1615207127_461;
   assign v3_1615207127_461 = v3_1615207127_49 ? v3_1615207127_470 : v3_1615207127_462;
   assign v3_1615207127_462 = v3_1615207127_46 ? v3_1615207127_469 : v3_1615207127_463;
   assign v3_1615207127_463 = v3_1615207127_43 ? v3_1615207127_465 : v3_1615207127_464;
   assign v3_1615207127_464 = v3_1615207127_23;
   assign v3_1615207127_465 = v3_1615207127_42 ? v3_1615207127_467 : v3_1615207127_466;
   assign v3_1615207127_466 = v3_1615207127_23;
   assign v3_1615207127_467 = v3_1615207127_468;
   assign v3_1615207127_468 = v3_1615207127_23 + v3_1615207127_10;
   assign v3_1615207127_469 = v3_1615207127_23;
   assign v3_1615207127_470 = v3_1615207127_23;
   assign v3_1615207127_471 = v3_1615207127_59 ? v3_1615207127_473 : v3_1615207127_472;
   assign v3_1615207127_472 = v3_1615207127_23;
   assign v3_1615207127_473 = v3_1615207127_58 ? v3_1615207127_476 : v3_1615207127_474;
   assign v3_1615207127_474 = v3_1615207127_475;
   assign v3_1615207127_475 = v3_1615207127_23 - v3_1615207127_55;
   assign v3_1615207127_476 = v3_1615207127_23;
   assign v3_1615207127_477 = v3_1615207127_23;
   assign v3_1615207127_478 = v3_1615207127_23;
   assign v3_1615207127_479 = v3_1615207127_70 ? v3_1615207127_481 : v3_1615207127_480;
   assign v3_1615207127_480 = v3_1615207127_23;
   assign v3_1615207127_481 = v3_1615207127_485 ? v3_1615207127_484 : v3_1615207127_482;
   assign v3_1615207127_482 = v3_1615207127_483;
   assign v3_1615207127_483 = v3_1615207127_23 + coinInA;
   assign v3_1615207127_484 = 6'b111111; 
   assign v3_1615207127_485 = v3_1615207127_486 >= v3_1615207127_492;
   assign v3_1615207127_486 = v3_1615207127_491;
   assign v3_1615207127_487 = v3_1615207127_488;
   assign v3_1615207127_488 = {v3_1615207127_252, v3_1615207127_23};
   assign v3_1615207127_489 = v3_1615207127_490;
   assign v3_1615207127_490 = {v3_1615207127_252, coinInA};
   assign v3_1615207127_491 = v3_1615207127_487 + v3_1615207127_489;
   assign v3_1615207127_492 = 7'b0111111; 
   assign v3_1615207127_493 = v3_1615207127_494;
   assign v3_1615207127_494 = 6'b000101; 
   assign v3_1615207127_495 = 6'b000000; 
   assign v3_1615207127_496 = v3_1615207127_75 ? v3_1615207127_533 : v3_1615207127_497;
   assign v3_1615207127_497 = v3_1615207127_17 ? v3_1615207127_499 : v3_1615207127_498;
   assign v3_1615207127_498 = v3_1615207127_24;
   assign v3_1615207127_499 = v3_1615207127_73 ? v3_1615207127_521 : v3_1615207127_500;
   assign v3_1615207127_500 = v3_1615207127_66 ? v3_1615207127_520 : v3_1615207127_501;
   assign v3_1615207127_501 = v3_1615207127_64 ? v3_1615207127_519 : v3_1615207127_502;
   assign v3_1615207127_502 = v3_1615207127_61 ? v3_1615207127_518 : v3_1615207127_503;
   assign v3_1615207127_503 = v3_1615207127_49 ? v3_1615207127_512 : v3_1615207127_504;
   assign v3_1615207127_504 = v3_1615207127_46 ? v3_1615207127_511 : v3_1615207127_505;
   assign v3_1615207127_505 = v3_1615207127_43 ? v3_1615207127_507 : v3_1615207127_506;
   assign v3_1615207127_506 = v3_1615207127_24;
   assign v3_1615207127_507 = v3_1615207127_42 ? v3_1615207127_509 : v3_1615207127_508;
   assign v3_1615207127_508 = v3_1615207127_24;
   assign v3_1615207127_509 = v3_1615207127_510;
   assign v3_1615207127_510 = v3_1615207127_24 + v3_1615207127_11;
   assign v3_1615207127_511 = v3_1615207127_24;
   assign v3_1615207127_512 = v3_1615207127_99 ? v3_1615207127_514 : v3_1615207127_513;
   assign v3_1615207127_513 = v3_1615207127_24;
   assign v3_1615207127_514 = v3_1615207127_98 ? v3_1615207127_517 : v3_1615207127_515;
   assign v3_1615207127_515 = v3_1615207127_516;
   assign v3_1615207127_516 = v3_1615207127_24 - v3_1615207127_55;
   assign v3_1615207127_517 = v3_1615207127_24;
   assign v3_1615207127_518 = v3_1615207127_24;
   assign v3_1615207127_519 = v3_1615207127_24;
   assign v3_1615207127_520 = v3_1615207127_24;
   assign v3_1615207127_521 = v3_1615207127_70 ? v3_1615207127_523 : v3_1615207127_522;
   assign v3_1615207127_522 = v3_1615207127_24;
   assign v3_1615207127_523 = v3_1615207127_526 ? v3_1615207127_484 : v3_1615207127_524;
   assign v3_1615207127_524 = v3_1615207127_525;
   assign v3_1615207127_525 = v3_1615207127_24 + coinInB;
   assign v3_1615207127_526 = v3_1615207127_527 >= v3_1615207127_492;
   assign v3_1615207127_527 = v3_1615207127_532;
   assign v3_1615207127_528 = v3_1615207127_529;
   assign v3_1615207127_529 = {v3_1615207127_252, v3_1615207127_24};
   assign v3_1615207127_530 = v3_1615207127_531;
   assign v3_1615207127_531 = {v3_1615207127_252, coinInB};
   assign v3_1615207127_532 = v3_1615207127_528 + v3_1615207127_530;
   assign v3_1615207127_533 = v3_1615207127_534;
   assign v3_1615207127_534 = 6'b011110; 
   assign v3_1615207127_535 = 6'b000000; 
   assign v3_1615207127_536 = v3_1615207127_75 ? v3_1615207127_569 : v3_1615207127_537;
   assign v3_1615207127_537 = v3_1615207127_17 ? v3_1615207127_539 : v3_1615207127_538;
   assign v3_1615207127_538 = v3_1615207127_25;
   assign v3_1615207127_539 = v3_1615207127_73 ? v3_1615207127_557 : v3_1615207127_540;
   assign v3_1615207127_540 = v3_1615207127_66 ? v3_1615207127_556 : v3_1615207127_541;
   assign v3_1615207127_541 = v3_1615207127_64 ? v3_1615207127_555 : v3_1615207127_542;
   assign v3_1615207127_542 = v3_1615207127_61 ? v3_1615207127_554 : v3_1615207127_543;
   assign v3_1615207127_543 = v3_1615207127_49 ? v3_1615207127_553 : v3_1615207127_544;
   assign v3_1615207127_544 = v3_1615207127_46 ? v3_1615207127_552 : v3_1615207127_545;
   assign v3_1615207127_545 = v3_1615207127_43 ? v3_1615207127_547 : v3_1615207127_546;
   assign v3_1615207127_546 = v3_1615207127_25;
   assign v3_1615207127_547 = v3_1615207127_42 ? v3_1615207127_550 : v3_1615207127_548;
   assign v3_1615207127_548 = v3_1615207127_549;
   assign v3_1615207127_549 = v3_1615207127_25 - v3_1615207127_55;
   assign v3_1615207127_550 = v3_1615207127_551;
   assign v3_1615207127_551 = v3_1615207127_25 + v3_1615207127_13;
   assign v3_1615207127_552 = v3_1615207127_25;
   assign v3_1615207127_553 = v3_1615207127_25;
   assign v3_1615207127_554 = v3_1615207127_25;
   assign v3_1615207127_555 = v3_1615207127_25;
   assign v3_1615207127_556 = v3_1615207127_25;
   assign v3_1615207127_557 = v3_1615207127_70 ? v3_1615207127_559 : v3_1615207127_558;
   assign v3_1615207127_558 = v3_1615207127_25;
   assign v3_1615207127_559 = v3_1615207127_562 ? v3_1615207127_484 : v3_1615207127_560;
   assign v3_1615207127_560 = v3_1615207127_561;
   assign v3_1615207127_561 = v3_1615207127_25 + coinInD;
   assign v3_1615207127_562 = v3_1615207127_563 >= v3_1615207127_492;
   assign v3_1615207127_563 = v3_1615207127_568;
   assign v3_1615207127_564 = v3_1615207127_565;
   assign v3_1615207127_565 = {v3_1615207127_252, v3_1615207127_25};
   assign v3_1615207127_566 = v3_1615207127_567;
   assign v3_1615207127_567 = {v3_1615207127_252, coinInD};
   assign v3_1615207127_568 = v3_1615207127_564 + v3_1615207127_566;
   assign v3_1615207127_569 = v3_1615207127_570;
   assign v3_1615207127_570 = 6'b010100; 
   assign v3_1615207127_571 = 6'b000000; 
   assign v3_1615207127_572 = v3_1615207127_75 ? v3_1615207127_609 : v3_1615207127_573;
   assign v3_1615207127_573 = v3_1615207127_17 ? v3_1615207127_575 : v3_1615207127_574;
   assign v3_1615207127_574 = v3_1615207127_26;
   assign v3_1615207127_575 = v3_1615207127_73 ? v3_1615207127_597 : v3_1615207127_576;
   assign v3_1615207127_576 = v3_1615207127_66 ? v3_1615207127_596 : v3_1615207127_577;
   assign v3_1615207127_577 = v3_1615207127_64 ? v3_1615207127_595 : v3_1615207127_578;
   assign v3_1615207127_578 = v3_1615207127_61 ? v3_1615207127_594 : v3_1615207127_579;
   assign v3_1615207127_579 = v3_1615207127_49 ? v3_1615207127_593 : v3_1615207127_580;
   assign v3_1615207127_580 = v3_1615207127_46 ? v3_1615207127_587 : v3_1615207127_581;
   assign v3_1615207127_581 = v3_1615207127_43 ? v3_1615207127_583 : v3_1615207127_582;
   assign v3_1615207127_582 = v3_1615207127_26;
   assign v3_1615207127_583 = v3_1615207127_42 ? v3_1615207127_585 : v3_1615207127_584;
   assign v3_1615207127_584 = v3_1615207127_26;
   assign v3_1615207127_585 = v3_1615207127_586;
   assign v3_1615207127_586 = v3_1615207127_26 + v3_1615207127_12;
   assign v3_1615207127_587 = v3_1615207127_130 ? v3_1615207127_589 : v3_1615207127_588;
   assign v3_1615207127_588 = v3_1615207127_26;
   assign v3_1615207127_589 = v3_1615207127_129 ? v3_1615207127_592 : v3_1615207127_590;
   assign v3_1615207127_590 = v3_1615207127_591;
   assign v3_1615207127_591 = v3_1615207127_26 - v3_1615207127_55;
   assign v3_1615207127_592 = v3_1615207127_26;
   assign v3_1615207127_593 = v3_1615207127_26;
   assign v3_1615207127_594 = v3_1615207127_26;
   assign v3_1615207127_595 = v3_1615207127_26;
   assign v3_1615207127_596 = v3_1615207127_26;
   assign v3_1615207127_597 = v3_1615207127_70 ? v3_1615207127_599 : v3_1615207127_598;
   assign v3_1615207127_598 = v3_1615207127_26;
   assign v3_1615207127_599 = v3_1615207127_602 ? v3_1615207127_484 : v3_1615207127_600;
   assign v3_1615207127_600 = v3_1615207127_601;
   assign v3_1615207127_601 = v3_1615207127_26 + coinInC;
   assign v3_1615207127_602 = v3_1615207127_603 >= v3_1615207127_492;
   assign v3_1615207127_603 = v3_1615207127_608;
   assign v3_1615207127_604 = v3_1615207127_605;
   assign v3_1615207127_605 = {v3_1615207127_252, v3_1615207127_26};
   assign v3_1615207127_606 = v3_1615207127_607;
   assign v3_1615207127_607 = {v3_1615207127_252, coinInC};
   assign v3_1615207127_608 = v3_1615207127_604 + v3_1615207127_606;
   assign v3_1615207127_609 = v3_1615207127_610;
   assign v3_1615207127_610 = 6'b001010; 
   assign v3_1615207127_611 = 6'b000000; 

   // Output Net Assignments
   assign coinOutA = v3_1615207127_10;
   assign coinOutB = v3_1615207127_11;
   assign coinOutC = v3_1615207127_12;
   assign coinOutD = v3_1615207127_13;
   assign itemTypeOut = v3_1615207127_14;
   assign itemNumberOut = v3_1615207127_15;
   assign serviceTypeOut = v3_1615207127_16;

   // Non-blocking Assignments
   always @ (posedge clk) begin
      v3_1615207127_10 <= v3_1615207127_27;
      v3_1615207127_11 <= v3_1615207127_77;
      v3_1615207127_12 <= v3_1615207127_109;
      v3_1615207127_13 <= v3_1615207127_141;
      v3_1615207127_14 <= v3_1615207127_166;
      v3_1615207127_15 <= v3_1615207127_176;
      v3_1615207127_16 <= v3_1615207127_209;
      v3_1615207127_17 <= v3_1615207127_231;
      v3_1615207127_18 <= v3_1615207127_236;
      v3_1615207127_19 <= v3_1615207127_255;
      v3_1615207127_20 <= v3_1615207127_292;
      v3_1615207127_21 <= v3_1615207127_302;
      v3_1615207127_22 <= v3_1615207127_335;
      v3_1615207127_23 <= v3_1615207127_454;
      v3_1615207127_24 <= v3_1615207127_496;
      v3_1615207127_25 <= v3_1615207127_536;
      v3_1615207127_26 <= v3_1615207127_572;
   end
endmodule
