// RTL (Verilog) generated @ Thu Jun  3 01:48:56 2021 by V3 
//               compiled @ Mar  8 2021 00:47:13
// Internal nets are renamed with prefix "v3_1622710136_".

// Module vendingMachine
module vendingMachine
(
   clk,
   reset,
   coinInNTD_50,
   coinInNTD_10,
   coinInNTD_5,
   coinInNTD_1,
   itemTypeIn,
   p,
   coinOutNTD_50,
   coinOutNTD_10,
   coinOutNTD_5,
   coinOutNTD_1,
   itemTypeOut,
   serviceTypeOut
);

   // Clock Signal for Synchronous DFF
   input clk;

   // I/O Declarations
   input reset;
   input [1:0] coinInNTD_50;
   input [1:0] coinInNTD_10;
   input [1:0] coinInNTD_5;
   input [1:0] coinInNTD_1;
   input [1:0] itemTypeIn;
   output p;
   output [2:0] coinOutNTD_50;
   output [2:0] coinOutNTD_10;
   output [2:0] coinOutNTD_5;
   output [2:0] coinOutNTD_1;
   output [1:0] itemTypeOut;
   output [1:0] serviceTypeOut;

   // Wire and Reg Declarations
   wire v3_1622710136_0;
   wire clk;
   wire reset;
   wire [1:0] coinInNTD_50;
   wire [1:0] coinInNTD_10;
   wire [1:0] coinInNTD_5;
   wire [1:0] coinInNTD_1;
   wire [1:0] itemTypeIn;
   reg [2:0] v3_1622710136_8;
   reg [2:0] v3_1622710136_9;
   reg [2:0] v3_1622710136_10;
   reg [2:0] v3_1622710136_11;
   reg [1:0] v3_1622710136_12;
   reg [1:0] v3_1622710136_13;
   reg v3_1622710136_14;
   reg [7:0] v3_1622710136_15;
   reg v3_1622710136_16;
   reg [1:0] v3_1622710136_17;
   reg [7:0] v3_1622710136_18;
   reg [2:0] v3_1622710136_19;
   reg [2:0] v3_1622710136_20;
   reg [2:0] v3_1622710136_21;
   reg [2:0] v3_1622710136_22;
   wire [2:0] v3_1622710136_23;
   wire [2:0] v3_1622710136_24;
   wire [2:0] v3_1622710136_25;
   wire [2:0] v3_1622710136_26;
   wire [2:0] v3_1622710136_27;
   wire [2:0] v3_1622710136_28;
   wire [2:0] v3_1622710136_29;
   wire [2:0] v3_1622710136_30;
   wire [2:0] v3_1622710136_31;
   wire [2:0] v3_1622710136_32;
   wire [2:0] v3_1622710136_33;
   wire [2:0] v3_1622710136_34;
   wire [2:0] v3_1622710136_35;
   wire v3_1622710136_36;
   wire v3_1622710136_37;
   wire [7:0] v3_1622710136_38;
   wire v3_1622710136_39;
   wire [1:0] v3_1622710136_40;
   wire v3_1622710136_41;
   wire [1:0] v3_1622710136_42;
   wire [2:0] v3_1622710136_43;
   wire [2:0] v3_1622710136_44;
   wire [2:0] v3_1622710136_45;
   wire [2:0] v3_1622710136_46;
   wire [2:0] v3_1622710136_47;
   wire v3_1622710136_48;
   wire v3_1622710136_49;
   wire [7:0] v3_1622710136_50;
   wire v3_1622710136_51;
   wire [1:0] v3_1622710136_52;
   wire v3_1622710136_53;
   wire [2:0] v3_1622710136_54;
   wire v3_1622710136_55;
   wire [2:0] v3_1622710136_56;
   wire [2:0] v3_1622710136_57;
   wire v3_1622710136_58;
   wire v3_1622710136_59;
   wire v3_1622710136_60;
   wire [2:0] v3_1622710136_61;
   wire v3_1622710136_62;
   wire [2:0] v3_1622710136_63;
   wire [2:0] v3_1622710136_64;
   wire [2:0] v3_1622710136_65;
   wire [2:0] v3_1622710136_66;
   wire [2:0] v3_1622710136_67;
   wire [2:0] v3_1622710136_68;
   wire [2:0] v3_1622710136_69;
   wire [2:0] v3_1622710136_70;
   wire [2:0] v3_1622710136_71;
   wire [2:0] v3_1622710136_72;
   wire [2:0] v3_1622710136_73;
   wire [2:0] v3_1622710136_74;
   wire [2:0] v3_1622710136_75;
   wire [2:0] v3_1622710136_76;
   wire [2:0] v3_1622710136_77;
   wire [2:0] v3_1622710136_78;
   wire [2:0] v3_1622710136_79;
   wire v3_1622710136_80;
   wire v3_1622710136_81;
   wire [7:0] v3_1622710136_82;
   wire [2:0] v3_1622710136_83;
   wire [2:0] v3_1622710136_84;
   wire [2:0] v3_1622710136_85;
   wire [2:0] v3_1622710136_86;
   wire [2:0] v3_1622710136_87;
   wire [2:0] v3_1622710136_88;
   wire [2:0] v3_1622710136_89;
   wire [2:0] v3_1622710136_90;
   wire [2:0] v3_1622710136_91;
   wire [2:0] v3_1622710136_92;
   wire [2:0] v3_1622710136_93;
   wire [2:0] v3_1622710136_94;
   wire [2:0] v3_1622710136_95;
   wire [2:0] v3_1622710136_96;
   wire [2:0] v3_1622710136_97;
   wire [2:0] v3_1622710136_98;
   wire [2:0] v3_1622710136_99;
   wire [2:0] v3_1622710136_100;
   wire [2:0] v3_1622710136_101;
   wire [2:0] v3_1622710136_102;
   wire [2:0] v3_1622710136_103;
   wire v3_1622710136_104;
   wire v3_1622710136_105;
   wire [7:0] v3_1622710136_106;
   wire [2:0] v3_1622710136_107;
   wire [2:0] v3_1622710136_108;
   wire [2:0] v3_1622710136_109;
   wire [2:0] v3_1622710136_110;
   wire [2:0] v3_1622710136_111;
   wire [2:0] v3_1622710136_112;
   wire [2:0] v3_1622710136_113;
   wire [2:0] v3_1622710136_114;
   wire [2:0] v3_1622710136_115;
   wire [2:0] v3_1622710136_116;
   wire [2:0] v3_1622710136_117;
   wire [2:0] v3_1622710136_118;
   wire [2:0] v3_1622710136_119;
   wire [2:0] v3_1622710136_120;
   wire [2:0] v3_1622710136_121;
   wire [2:0] v3_1622710136_122;
   wire [2:0] v3_1622710136_123;
   wire [2:0] v3_1622710136_124;
   wire [2:0] v3_1622710136_125;
   wire [2:0] v3_1622710136_126;
   wire [2:0] v3_1622710136_127;
   wire [2:0] v3_1622710136_128;
   wire [2:0] v3_1622710136_129;
   wire [2:0] v3_1622710136_130;
   wire [1:0] v3_1622710136_131;
   wire [1:0] v3_1622710136_132;
   wire [1:0] v3_1622710136_133;
   wire [1:0] v3_1622710136_134;
   wire [1:0] v3_1622710136_135;
   wire [1:0] v3_1622710136_136;
   wire [1:0] v3_1622710136_137;
   wire [1:0] v3_1622710136_138;
   wire [1:0] v3_1622710136_139;
   wire [1:0] v3_1622710136_140;
   wire [1:0] v3_1622710136_141;
   wire [1:0] v3_1622710136_142;
   wire [1:0] v3_1622710136_143;
   wire [1:0] v3_1622710136_144;
   wire v3_1622710136_145;
   wire v3_1622710136_146;
   wire [1:0] v3_1622710136_147;
   wire [1:0] v3_1622710136_148;
   wire [1:0] v3_1622710136_149;
   wire [1:0] v3_1622710136_150;
   wire [1:0] v3_1622710136_151;
   wire [1:0] v3_1622710136_152;
   wire [1:0] v3_1622710136_153;
   wire [1:0] v3_1622710136_154;
   wire [1:0] v3_1622710136_155;
   wire [1:0] v3_1622710136_156;
   wire [1:0] v3_1622710136_157;
   wire [1:0] v3_1622710136_158;
   wire [1:0] v3_1622710136_159;
   wire [1:0] v3_1622710136_160;
   wire [1:0] v3_1622710136_161;
   wire [1:0] v3_1622710136_162;
   wire [1:0] v3_1622710136_163;
   wire [1:0] v3_1622710136_164;
   wire [1:0] v3_1622710136_165;
   wire [1:0] v3_1622710136_166;
   wire [1:0] v3_1622710136_167;
   wire [1:0] v3_1622710136_168;
   wire [1:0] v3_1622710136_169;
   wire v3_1622710136_170;
   wire v3_1622710136_171;
   wire v3_1622710136_172;
   wire v3_1622710136_173;
   wire v3_1622710136_174;
   wire [7:0] v3_1622710136_175;
   wire [7:0] v3_1622710136_176;
   wire [7:0] v3_1622710136_177;
   wire [7:0] v3_1622710136_178;
   wire [7:0] v3_1622710136_179;
   wire [7:0] v3_1622710136_180;
   wire [7:0] v3_1622710136_181;
   wire [7:0] v3_1622710136_182;
   wire [7:0] v3_1622710136_183;
   wire [7:0] v3_1622710136_184;
   wire [5:0] v3_1622710136_185;
   wire [7:0] v3_1622710136_186;
   wire [7:0] v3_1622710136_187;
   wire [7:0] v3_1622710136_188;
   wire [7:0] v3_1622710136_189;
   wire [7:0] v3_1622710136_190;
   wire [7:0] v3_1622710136_191;
   wire [7:0] v3_1622710136_192;
   wire [7:0] v3_1622710136_193;
   wire [7:0] v3_1622710136_194;
   wire [7:0] v3_1622710136_195;
   wire [7:0] v3_1622710136_196;
   wire [7:0] v3_1622710136_197;
   wire [7:0] v3_1622710136_198;
   wire [7:0] v3_1622710136_199;
   wire [7:0] v3_1622710136_200;
   wire [7:0] v3_1622710136_201;
   wire [7:0] v3_1622710136_202;
   wire [7:0] v3_1622710136_203;
   wire [7:0] v3_1622710136_204;
   wire [7:0] v3_1622710136_205;
   wire v3_1622710136_206;
   wire v3_1622710136_207;
   wire v3_1622710136_208;
   wire v3_1622710136_209;
   wire v3_1622710136_210;
   wire v3_1622710136_211;
   wire v3_1622710136_212;
   wire v3_1622710136_213;
   wire v3_1622710136_214;
   wire v3_1622710136_215;
   wire v3_1622710136_216;
   wire v3_1622710136_217;
   wire v3_1622710136_218;
   wire v3_1622710136_219;
   wire [1:0] v3_1622710136_220;
   wire [1:0] v3_1622710136_221;
   wire [1:0] v3_1622710136_222;
   wire [1:0] v3_1622710136_223;
   wire [1:0] v3_1622710136_224;
   wire [1:0] v3_1622710136_225;
   wire [1:0] v3_1622710136_226;
   wire [1:0] v3_1622710136_227;
   wire [1:0] v3_1622710136_228;
   wire [1:0] v3_1622710136_229;
   wire [1:0] v3_1622710136_230;
   wire [1:0] v3_1622710136_231;
   wire [1:0] v3_1622710136_232;
   wire [1:0] v3_1622710136_233;
   wire [1:0] v3_1622710136_234;
   wire [1:0] v3_1622710136_235;
   wire [1:0] v3_1622710136_236;
   wire [1:0] v3_1622710136_237;
   wire [1:0] v3_1622710136_238;
   wire [1:0] v3_1622710136_239;
   wire [1:0] v3_1622710136_240;
   wire [1:0] v3_1622710136_241;
   wire [1:0] v3_1622710136_242;
   wire [1:0] v3_1622710136_243;
   wire [1:0] v3_1622710136_244;
   wire [1:0] v3_1622710136_245;
   wire [1:0] v3_1622710136_246;
   wire [1:0] v3_1622710136_247;
   wire [1:0] v3_1622710136_248;
   wire [7:0] v3_1622710136_249;
   wire [7:0] v3_1622710136_250;
   wire [7:0] v3_1622710136_251;
   wire [7:0] v3_1622710136_252;
   wire [7:0] v3_1622710136_253;
   wire [7:0] v3_1622710136_254;
   wire [7:0] v3_1622710136_255;
   wire [7:0] v3_1622710136_256;
   wire [7:0] v3_1622710136_257;
   wire [7:0] v3_1622710136_258;
   wire [7:0] v3_1622710136_259;
   wire [7:0] v3_1622710136_260;
   wire [7:0] v3_1622710136_261;
   wire [7:0] v3_1622710136_262;
   wire [7:0] v3_1622710136_263;
   wire [7:0] v3_1622710136_264;
   wire [7:0] v3_1622710136_265;
   wire [7:0] v3_1622710136_266;
   wire [7:0] v3_1622710136_267;
   wire [7:0] v3_1622710136_268;
   wire [7:0] v3_1622710136_269;
   wire [7:0] v3_1622710136_270;
   wire [7:0] v3_1622710136_271;
   wire [7:0] v3_1622710136_272;
   wire [7:0] v3_1622710136_273;
   wire [7:0] v3_1622710136_274;
   wire [7:0] v3_1622710136_275;
   wire [7:0] v3_1622710136_276;
   wire [7:0] v3_1622710136_277;
   wire [7:0] v3_1622710136_278;
   wire [7:0] v3_1622710136_279;
   wire [7:0] v3_1622710136_280;
   wire [7:0] v3_1622710136_281;
   wire [7:0] v3_1622710136_282;
   wire [7:0] v3_1622710136_283;
   wire v3_1622710136_284;
   wire [7:0] v3_1622710136_285;
   wire v3_1622710136_286;
   wire [7:0] v3_1622710136_287;
   wire v3_1622710136_288;
   wire [7:0] v3_1622710136_289;
   wire [7:0] v3_1622710136_290;
   wire [2:0] v3_1622710136_291;
   wire [2:0] v3_1622710136_292;
   wire [2:0] v3_1622710136_293;
   wire [2:0] v3_1622710136_294;
   wire [2:0] v3_1622710136_295;
   wire [2:0] v3_1622710136_296;
   wire [2:0] v3_1622710136_297;
   wire [2:0] v3_1622710136_298;
   wire [2:0] v3_1622710136_299;
   wire [2:0] v3_1622710136_300;
   wire [2:0] v3_1622710136_301;
   wire [2:0] v3_1622710136_302;
   wire [2:0] v3_1622710136_303;
   wire [2:0] v3_1622710136_304;
   wire [2:0] v3_1622710136_305;
   wire [2:0] v3_1622710136_306;
   wire [2:0] v3_1622710136_307;
   wire [2:0] v3_1622710136_308;
   wire [2:0] v3_1622710136_309;
   wire [2:0] v3_1622710136_310;
   wire [2:0] v3_1622710136_311;
   wire [2:0] v3_1622710136_312;
   wire [2:0] v3_1622710136_313;
   wire [2:0] v3_1622710136_314;
   wire v3_1622710136_315;
   wire [3:0] v3_1622710136_316;
   wire [3:0] v3_1622710136_317;
   wire [3:0] v3_1622710136_318;
   wire [3:0] v3_1622710136_319;
   wire [3:0] v3_1622710136_320;
   wire [3:0] v3_1622710136_321;
   wire [3:0] v3_1622710136_322;
   wire [2:0] v3_1622710136_323;
   wire [2:0] v3_1622710136_324;
   wire [2:0] v3_1622710136_325;
   wire [2:0] v3_1622710136_326;
   wire [2:0] v3_1622710136_327;
   wire [2:0] v3_1622710136_328;
   wire [2:0] v3_1622710136_329;
   wire [2:0] v3_1622710136_330;
   wire [2:0] v3_1622710136_331;
   wire [2:0] v3_1622710136_332;
   wire [2:0] v3_1622710136_333;
   wire [2:0] v3_1622710136_334;
   wire [2:0] v3_1622710136_335;
   wire [2:0] v3_1622710136_336;
   wire [2:0] v3_1622710136_337;
   wire [2:0] v3_1622710136_338;
   wire [2:0] v3_1622710136_339;
   wire [2:0] v3_1622710136_340;
   wire [2:0] v3_1622710136_341;
   wire [2:0] v3_1622710136_342;
   wire [2:0] v3_1622710136_343;
   wire [2:0] v3_1622710136_344;
   wire [2:0] v3_1622710136_345;
   wire [2:0] v3_1622710136_346;
   wire [2:0] v3_1622710136_347;
   wire [2:0] v3_1622710136_348;
   wire v3_1622710136_349;
   wire [3:0] v3_1622710136_350;
   wire [3:0] v3_1622710136_351;
   wire [3:0] v3_1622710136_352;
   wire [3:0] v3_1622710136_353;
   wire [3:0] v3_1622710136_354;
   wire [3:0] v3_1622710136_355;
   wire [2:0] v3_1622710136_356;
   wire [2:0] v3_1622710136_357;
   wire [2:0] v3_1622710136_358;
   wire [2:0] v3_1622710136_359;
   wire [2:0] v3_1622710136_360;
   wire [2:0] v3_1622710136_361;
   wire [2:0] v3_1622710136_362;
   wire [2:0] v3_1622710136_363;
   wire [2:0] v3_1622710136_364;
   wire [2:0] v3_1622710136_365;
   wire [2:0] v3_1622710136_366;
   wire [2:0] v3_1622710136_367;
   wire [2:0] v3_1622710136_368;
   wire [2:0] v3_1622710136_369;
   wire [2:0] v3_1622710136_370;
   wire [2:0] v3_1622710136_371;
   wire [2:0] v3_1622710136_372;
   wire [2:0] v3_1622710136_373;
   wire [2:0] v3_1622710136_374;
   wire [2:0] v3_1622710136_375;
   wire [2:0] v3_1622710136_376;
   wire [2:0] v3_1622710136_377;
   wire [2:0] v3_1622710136_378;
   wire v3_1622710136_379;
   wire [3:0] v3_1622710136_380;
   wire [3:0] v3_1622710136_381;
   wire [3:0] v3_1622710136_382;
   wire [3:0] v3_1622710136_383;
   wire [3:0] v3_1622710136_384;
   wire [3:0] v3_1622710136_385;
   wire [2:0] v3_1622710136_386;
   wire [2:0] v3_1622710136_387;
   wire [2:0] v3_1622710136_388;
   wire [2:0] v3_1622710136_389;
   wire [2:0] v3_1622710136_390;
   wire [2:0] v3_1622710136_391;
   wire [2:0] v3_1622710136_392;
   wire [2:0] v3_1622710136_393;
   wire [2:0] v3_1622710136_394;
   wire [2:0] v3_1622710136_395;
   wire [2:0] v3_1622710136_396;
   wire [2:0] v3_1622710136_397;
   wire [2:0] v3_1622710136_398;
   wire [2:0] v3_1622710136_399;
   wire [2:0] v3_1622710136_400;
   wire [2:0] v3_1622710136_401;
   wire [2:0] v3_1622710136_402;
   wire [2:0] v3_1622710136_403;
   wire [2:0] v3_1622710136_404;
   wire [2:0] v3_1622710136_405;
   wire [2:0] v3_1622710136_406;
   wire [2:0] v3_1622710136_407;
   wire [2:0] v3_1622710136_408;
   wire [2:0] v3_1622710136_409;
   wire [2:0] v3_1622710136_410;
   wire v3_1622710136_411;
   wire [3:0] v3_1622710136_412;
   wire [3:0] v3_1622710136_413;
   wire [3:0] v3_1622710136_414;
   wire [3:0] v3_1622710136_415;
   wire [3:0] v3_1622710136_416;
   wire [3:0] v3_1622710136_417;
   wire [2:0] v3_1622710136_418;
   wire [2:0] v3_1622710136_419;
   wire v3_1622710136_420;
   wire v3_1622710136_421;
   wire v3_1622710136_422;
   wire v3_1622710136_423;
   wire v3_1622710136_424;
   wire v3_1622710136_425;
   wire v3_1622710136_426;
   wire v3_1622710136_427;
   wire [7:0] v3_1622710136_428;
   wire [7:0] v3_1622710136_429;
   wire [7:0] v3_1622710136_430;
   wire [7:0] v3_1622710136_431;
   wire [7:0] v3_1622710136_432;
   wire [4:0] v3_1622710136_433;
   wire [7:0] v3_1622710136_434;
   wire [7:0] v3_1622710136_435;
   wire [7:0] v3_1622710136_436;
   wire [7:0] v3_1622710136_437;
   wire [7:0] v3_1622710136_438;
   wire [7:0] v3_1622710136_439;
   wire [7:0] v3_1622710136_440;
   wire [7:0] v3_1622710136_441;
   wire [7:0] v3_1622710136_442;
   wire [7:0] v3_1622710136_443;
   wire [7:0] v3_1622710136_444;
   wire [7:0] v3_1622710136_445;
   wire [7:0] v3_1622710136_446;
   wire [7:0] v3_1622710136_447;
   wire [7:0] v3_1622710136_448;
   wire [7:0] v3_1622710136_449;
   wire [7:0] v3_1622710136_450;
   wire v3_1622710136_451;

   // Output Net Declarations
   wire p;
   wire [2:0] coinOutNTD_50;
   wire [2:0] coinOutNTD_10;
   wire [2:0] coinOutNTD_5;
   wire [2:0] coinOutNTD_1;
   wire [1:0] itemTypeOut;
   wire [1:0] serviceTypeOut;

   // Combinational Assignments
   assign v3_1622710136_0 = 1'b0; 
   assign v3_1622710136_23 = v3_1622710136_62 ? v3_1622710136_61 : v3_1622710136_24;
   assign v3_1622710136_24 = v3_1622710136_25;
   assign v3_1622710136_25 = v3_1622710136_60 ? v3_1622710136_56 : v3_1622710136_26;
   assign v3_1622710136_26 = v3_1622710136_55 ? v3_1622710136_54 : v3_1622710136_27;
   assign v3_1622710136_27 = v3_1622710136_53 ? v3_1622710136_32 : v3_1622710136_28;
   assign v3_1622710136_28 = v3_1622710136_51 ? v3_1622710136_43 : v3_1622710136_29;
   assign v3_1622710136_29 = v3_1622710136_41 ? v3_1622710136_32 : v3_1622710136_30;
   assign v3_1622710136_30 = v3_1622710136_39 ? v3_1622710136_32 : v3_1622710136_31;
   assign v3_1622710136_31 = v3_1622710136_37 ? v3_1622710136_33 : v3_1622710136_32;
   assign v3_1622710136_32 = v3_1622710136_8;
   assign v3_1622710136_33 = v3_1622710136_36 ? v3_1622710136_34 : v3_1622710136_32;
   assign v3_1622710136_34 = v3_1622710136_35;
   assign v3_1622710136_35 = 3'b000; 
   assign v3_1622710136_36 = v3_1622710136_21 == v3_1622710136_35;
   assign v3_1622710136_37 = v3_1622710136_18 >= v3_1622710136_38;
   assign v3_1622710136_38 = 8'b00000001; 
   assign v3_1622710136_39 = v3_1622710136_17 == v3_1622710136_40;
   assign v3_1622710136_40 = 2'b10; 
   assign v3_1622710136_41 = v3_1622710136_17 == v3_1622710136_42;
   assign v3_1622710136_42 = 2'b01; 
   assign v3_1622710136_43 = v3_1622710136_49 ? v3_1622710136_44 : v3_1622710136_32;
   assign v3_1622710136_44 = v3_1622710136_48 ? v3_1622710136_32 : v3_1622710136_45;
   assign v3_1622710136_45 = v3_1622710136_47;
   assign v3_1622710136_46 = 3'b001; 
   assign v3_1622710136_47 = v3_1622710136_8 + v3_1622710136_46;
   assign v3_1622710136_48 = v3_1622710136_19 == v3_1622710136_35;
   assign v3_1622710136_49 = v3_1622710136_18 >= v3_1622710136_50;
   assign v3_1622710136_50 = 8'b00110010; 
   assign v3_1622710136_51 = v3_1622710136_17 == v3_1622710136_52;
   assign v3_1622710136_52 = 2'b00; 
   assign v3_1622710136_53 = ~v3_1622710136_16;
   assign v3_1622710136_54 = v3_1622710136_35;
   assign v3_1622710136_55 = v3_1622710136_13 == v3_1622710136_52;
   assign v3_1622710136_56 = v3_1622710136_58 ? v3_1622710136_57 : v3_1622710136_32;
   assign v3_1622710136_57 = v3_1622710136_35;
   assign v3_1622710136_58 = ~v3_1622710136_59;
   assign v3_1622710136_59 = itemTypeIn == v3_1622710136_52;
   assign v3_1622710136_60 = v3_1622710136_13 == v3_1622710136_42;
   assign v3_1622710136_61 = v3_1622710136_35;
   assign v3_1622710136_62 = ~reset;
   assign v3_1622710136_63 = 3'b000; 
   assign v3_1622710136_64 = v3_1622710136_62 ? v3_1622710136_86 : v3_1622710136_65;
   assign v3_1622710136_65 = v3_1622710136_66;
   assign v3_1622710136_66 = v3_1622710136_60 ? v3_1622710136_84 : v3_1622710136_67;
   assign v3_1622710136_67 = v3_1622710136_55 ? v3_1622710136_83 : v3_1622710136_68;
   assign v3_1622710136_68 = v3_1622710136_53 ? v3_1622710136_73 : v3_1622710136_69;
   assign v3_1622710136_69 = v3_1622710136_51 ? v3_1622710136_73 : v3_1622710136_70;
   assign v3_1622710136_70 = v3_1622710136_41 ? v3_1622710136_76 : v3_1622710136_71;
   assign v3_1622710136_71 = v3_1622710136_39 ? v3_1622710136_73 : v3_1622710136_72;
   assign v3_1622710136_72 = v3_1622710136_37 ? v3_1622710136_74 : v3_1622710136_73;
   assign v3_1622710136_73 = v3_1622710136_9;
   assign v3_1622710136_74 = v3_1622710136_36 ? v3_1622710136_75 : v3_1622710136_73;
   assign v3_1622710136_75 = v3_1622710136_35;
   assign v3_1622710136_76 = v3_1622710136_81 ? v3_1622710136_77 : v3_1622710136_73;
   assign v3_1622710136_77 = v3_1622710136_80 ? v3_1622710136_73 : v3_1622710136_78;
   assign v3_1622710136_78 = v3_1622710136_79;
   assign v3_1622710136_79 = v3_1622710136_9 + v3_1622710136_46;
   assign v3_1622710136_80 = v3_1622710136_20 == v3_1622710136_35;
   assign v3_1622710136_81 = v3_1622710136_18 >= v3_1622710136_82;
   assign v3_1622710136_82 = 8'b00001010; 
   assign v3_1622710136_83 = v3_1622710136_35;
   assign v3_1622710136_84 = v3_1622710136_58 ? v3_1622710136_85 : v3_1622710136_73;
   assign v3_1622710136_85 = v3_1622710136_35;
   assign v3_1622710136_86 = v3_1622710136_35;
   assign v3_1622710136_87 = 3'b000; 
   assign v3_1622710136_88 = v3_1622710136_62 ? v3_1622710136_110 : v3_1622710136_89;
   assign v3_1622710136_89 = v3_1622710136_90;
   assign v3_1622710136_90 = v3_1622710136_60 ? v3_1622710136_108 : v3_1622710136_91;
   assign v3_1622710136_91 = v3_1622710136_55 ? v3_1622710136_107 : v3_1622710136_92;
   assign v3_1622710136_92 = v3_1622710136_53 ? v3_1622710136_97 : v3_1622710136_93;
   assign v3_1622710136_93 = v3_1622710136_51 ? v3_1622710136_97 : v3_1622710136_94;
   assign v3_1622710136_94 = v3_1622710136_41 ? v3_1622710136_97 : v3_1622710136_95;
   assign v3_1622710136_95 = v3_1622710136_39 ? v3_1622710136_100 : v3_1622710136_96;
   assign v3_1622710136_96 = v3_1622710136_37 ? v3_1622710136_98 : v3_1622710136_97;
   assign v3_1622710136_97 = v3_1622710136_10;
   assign v3_1622710136_98 = v3_1622710136_36 ? v3_1622710136_99 : v3_1622710136_97;
   assign v3_1622710136_99 = v3_1622710136_35;
   assign v3_1622710136_100 = v3_1622710136_105 ? v3_1622710136_101 : v3_1622710136_97;
   assign v3_1622710136_101 = v3_1622710136_104 ? v3_1622710136_97 : v3_1622710136_102;
   assign v3_1622710136_102 = v3_1622710136_103;
   assign v3_1622710136_103 = v3_1622710136_10 + v3_1622710136_46;
   assign v3_1622710136_104 = v3_1622710136_22 == v3_1622710136_35;
   assign v3_1622710136_105 = v3_1622710136_18 >= v3_1622710136_106;
   assign v3_1622710136_106 = 8'b00000101; 
   assign v3_1622710136_107 = v3_1622710136_35;
   assign v3_1622710136_108 = v3_1622710136_58 ? v3_1622710136_109 : v3_1622710136_97;
   assign v3_1622710136_109 = v3_1622710136_35;
   assign v3_1622710136_110 = v3_1622710136_35;
   assign v3_1622710136_111 = 3'b000; 
   assign v3_1622710136_112 = v3_1622710136_62 ? v3_1622710136_129 : v3_1622710136_113;
   assign v3_1622710136_113 = v3_1622710136_114;
   assign v3_1622710136_114 = v3_1622710136_60 ? v3_1622710136_127 : v3_1622710136_115;
   assign v3_1622710136_115 = v3_1622710136_55 ? v3_1622710136_126 : v3_1622710136_116;
   assign v3_1622710136_116 = v3_1622710136_53 ? v3_1622710136_121 : v3_1622710136_117;
   assign v3_1622710136_117 = v3_1622710136_51 ? v3_1622710136_121 : v3_1622710136_118;
   assign v3_1622710136_118 = v3_1622710136_41 ? v3_1622710136_121 : v3_1622710136_119;
   assign v3_1622710136_119 = v3_1622710136_39 ? v3_1622710136_121 : v3_1622710136_120;
   assign v3_1622710136_120 = v3_1622710136_37 ? v3_1622710136_122 : v3_1622710136_121;
   assign v3_1622710136_121 = v3_1622710136_11;
   assign v3_1622710136_122 = v3_1622710136_36 ? v3_1622710136_125 : v3_1622710136_123;
   assign v3_1622710136_123 = v3_1622710136_124;
   assign v3_1622710136_124 = v3_1622710136_11 + v3_1622710136_46;
   assign v3_1622710136_125 = v3_1622710136_35;
   assign v3_1622710136_126 = v3_1622710136_35;
   assign v3_1622710136_127 = v3_1622710136_58 ? v3_1622710136_128 : v3_1622710136_121;
   assign v3_1622710136_128 = v3_1622710136_35;
   assign v3_1622710136_129 = v3_1622710136_35;
   assign v3_1622710136_130 = 3'b000; 
   assign v3_1622710136_131 = v3_1622710136_62 ? v3_1622710136_150 : v3_1622710136_132;
   assign v3_1622710136_132 = v3_1622710136_133;
   assign v3_1622710136_133 = v3_1622710136_60 ? v3_1622710136_148 : v3_1622710136_134;
   assign v3_1622710136_134 = v3_1622710136_55 ? v3_1622710136_147 : v3_1622710136_135;
   assign v3_1622710136_135 = v3_1622710136_53 ? v3_1622710136_143 : v3_1622710136_136;
   assign v3_1622710136_136 = v3_1622710136_51 ? v3_1622710136_140 : v3_1622710136_137;
   assign v3_1622710136_137 = v3_1622710136_41 ? v3_1622710136_140 : v3_1622710136_138;
   assign v3_1622710136_138 = v3_1622710136_39 ? v3_1622710136_140 : v3_1622710136_139;
   assign v3_1622710136_139 = v3_1622710136_37 ? v3_1622710136_141 : v3_1622710136_140;
   assign v3_1622710136_140 = v3_1622710136_12;
   assign v3_1622710136_141 = v3_1622710136_36 ? v3_1622710136_142 : v3_1622710136_140;
   assign v3_1622710136_142 = v3_1622710136_52;
   assign v3_1622710136_143 = v3_1622710136_145 ? v3_1622710136_144 : v3_1622710136_140;
   assign v3_1622710136_144 = v3_1622710136_52;
   assign v3_1622710136_145 = ~v3_1622710136_146;
   assign v3_1622710136_146 = v3_1622710136_15 >= v3_1622710136_18;
   assign v3_1622710136_147 = v3_1622710136_52;
   assign v3_1622710136_148 = v3_1622710136_58 ? v3_1622710136_149 : v3_1622710136_140;
   assign v3_1622710136_149 = itemTypeIn;
   assign v3_1622710136_150 = v3_1622710136_52;
   assign v3_1622710136_151 = 2'b00; 
   assign v3_1622710136_152 = v3_1622710136_62 ? v3_1622710136_168 : v3_1622710136_153;
   assign v3_1622710136_153 = v3_1622710136_154;
   assign v3_1622710136_154 = v3_1622710136_60 ? v3_1622710136_166 : v3_1622710136_155;
   assign v3_1622710136_155 = v3_1622710136_55 ? v3_1622710136_165 : v3_1622710136_156;
   assign v3_1622710136_156 = v3_1622710136_53 ? v3_1622710136_163 : v3_1622710136_157;
   assign v3_1622710136_157 = v3_1622710136_51 ? v3_1622710136_163 : v3_1622710136_158;
   assign v3_1622710136_158 = v3_1622710136_41 ? v3_1622710136_163 : v3_1622710136_159;
   assign v3_1622710136_159 = v3_1622710136_39 ? v3_1622710136_163 : v3_1622710136_160;
   assign v3_1622710136_160 = v3_1622710136_37 ? v3_1622710136_162 : v3_1622710136_161;
   assign v3_1622710136_161 = v3_1622710136_52;
   assign v3_1622710136_162 = v3_1622710136_36 ? v3_1622710136_164 : v3_1622710136_163;
   assign v3_1622710136_163 = v3_1622710136_13;
   assign v3_1622710136_164 = v3_1622710136_52;
   assign v3_1622710136_165 = v3_1622710136_42;
   assign v3_1622710136_166 = v3_1622710136_58 ? v3_1622710136_167 : v3_1622710136_163;
   assign v3_1622710136_167 = v3_1622710136_40;
   assign v3_1622710136_168 = v3_1622710136_42;
   assign v3_1622710136_169 = 2'b00; 
   assign v3_1622710136_170 = v3_1622710136_62 ? v3_1622710136_172 : v3_1622710136_171;
   assign v3_1622710136_171 = v3_1622710136_14;
   assign v3_1622710136_172 = v3_1622710136_173;
   assign v3_1622710136_173 = 1'b1; 
   assign v3_1622710136_174 = 1'b0; 
   assign v3_1622710136_175 = v3_1622710136_62 ? v3_1622710136_203 : v3_1622710136_176;
   assign v3_1622710136_176 = v3_1622710136_177;
   assign v3_1622710136_177 = v3_1622710136_60 ? v3_1622710136_179 : v3_1622710136_178;
   assign v3_1622710136_178 = v3_1622710136_15;
   assign v3_1622710136_179 = v3_1622710136_58 ? v3_1622710136_180 : v3_1622710136_178;
   assign v3_1622710136_180 = v3_1622710136_202;
   assign v3_1622710136_181 = v3_1622710136_197;
   assign v3_1622710136_182 = v3_1622710136_192;
   assign v3_1622710136_183 = v3_1622710136_187;
   assign v3_1622710136_184 = v3_1622710136_186;
   assign v3_1622710136_185 = 6'b000000; 
   assign v3_1622710136_186 = {v3_1622710136_185, coinInNTD_50};
   assign v3_1622710136_187 = v3_1622710136_50 * v3_1622710136_184;
   assign v3_1622710136_188 = v3_1622710136_191;
   assign v3_1622710136_189 = v3_1622710136_190;
   assign v3_1622710136_190 = {v3_1622710136_185, coinInNTD_10};
   assign v3_1622710136_191 = v3_1622710136_82 * v3_1622710136_189;
   assign v3_1622710136_192 = v3_1622710136_183 + v3_1622710136_188;
   assign v3_1622710136_193 = v3_1622710136_196;
   assign v3_1622710136_194 = v3_1622710136_195;
   assign v3_1622710136_195 = {v3_1622710136_185, coinInNTD_5};
   assign v3_1622710136_196 = v3_1622710136_106 * v3_1622710136_194;
   assign v3_1622710136_197 = v3_1622710136_182 + v3_1622710136_193;
   assign v3_1622710136_198 = v3_1622710136_201;
   assign v3_1622710136_199 = v3_1622710136_200;
   assign v3_1622710136_200 = {v3_1622710136_185, coinInNTD_1};
   assign v3_1622710136_201 = v3_1622710136_38 * v3_1622710136_199;
   assign v3_1622710136_202 = v3_1622710136_181 + v3_1622710136_198;
   assign v3_1622710136_203 = v3_1622710136_204;
   assign v3_1622710136_204 = 8'b00000000; 
   assign v3_1622710136_205 = 8'b00000000; 
   assign v3_1622710136_206 = v3_1622710136_62 ? v3_1622710136_218 : v3_1622710136_207;
   assign v3_1622710136_207 = v3_1622710136_208;
   assign v3_1622710136_208 = v3_1622710136_60 ? v3_1622710136_215 : v3_1622710136_209;
   assign v3_1622710136_209 = v3_1622710136_55 ? v3_1622710136_211 : v3_1622710136_210;
   assign v3_1622710136_210 = v3_1622710136_53 ? v3_1622710136_212 : v3_1622710136_211;
   assign v3_1622710136_211 = v3_1622710136_16;
   assign v3_1622710136_212 = v3_1622710136_145 ? v3_1622710136_214 : v3_1622710136_213;
   assign v3_1622710136_213 = v3_1622710136_173;
   assign v3_1622710136_214 = v3_1622710136_173;
   assign v3_1622710136_215 = v3_1622710136_58 ? v3_1622710136_216 : v3_1622710136_211;
   assign v3_1622710136_216 = v3_1622710136_217;
   assign v3_1622710136_217 = 1'b0; 
   assign v3_1622710136_218 = v3_1622710136_217;
   assign v3_1622710136_219 = 1'b0; 
   assign v3_1622710136_220 = v3_1622710136_62 ? v3_1622710136_247 : v3_1622710136_221;
   assign v3_1622710136_221 = v3_1622710136_222;
   assign v3_1622710136_222 = v3_1622710136_60 ? v3_1622710136_245 : v3_1622710136_223;
   assign v3_1622710136_223 = v3_1622710136_55 ? v3_1622710136_229 : v3_1622710136_224;
   assign v3_1622710136_224 = v3_1622710136_53 ? v3_1622710136_229 : v3_1622710136_225;
   assign v3_1622710136_225 = v3_1622710136_51 ? v3_1622710136_241 : v3_1622710136_226;
   assign v3_1622710136_226 = v3_1622710136_41 ? v3_1622710136_237 : v3_1622710136_227;
   assign v3_1622710136_227 = v3_1622710136_39 ? v3_1622710136_232 : v3_1622710136_228;
   assign v3_1622710136_228 = v3_1622710136_37 ? v3_1622710136_230 : v3_1622710136_229;
   assign v3_1622710136_229 = v3_1622710136_17;
   assign v3_1622710136_230 = v3_1622710136_36 ? v3_1622710136_231 : v3_1622710136_229;
   assign v3_1622710136_231 = v3_1622710136_52;
   assign v3_1622710136_232 = v3_1622710136_105 ? v3_1622710136_235 : v3_1622710136_233;
   assign v3_1622710136_233 = v3_1622710136_234;
   assign v3_1622710136_234 = 2'b11; 
   assign v3_1622710136_235 = v3_1622710136_104 ? v3_1622710136_236 : v3_1622710136_229;
   assign v3_1622710136_236 = v3_1622710136_234;
   assign v3_1622710136_237 = v3_1622710136_81 ? v3_1622710136_239 : v3_1622710136_238;
   assign v3_1622710136_238 = v3_1622710136_40;
   assign v3_1622710136_239 = v3_1622710136_80 ? v3_1622710136_240 : v3_1622710136_229;
   assign v3_1622710136_240 = v3_1622710136_40;
   assign v3_1622710136_241 = v3_1622710136_49 ? v3_1622710136_243 : v3_1622710136_242;
   assign v3_1622710136_242 = v3_1622710136_42;
   assign v3_1622710136_243 = v3_1622710136_48 ? v3_1622710136_244 : v3_1622710136_229;
   assign v3_1622710136_244 = v3_1622710136_42;
   assign v3_1622710136_245 = v3_1622710136_58 ? v3_1622710136_246 : v3_1622710136_229;
   assign v3_1622710136_246 = v3_1622710136_52;
   assign v3_1622710136_247 = v3_1622710136_52;
   assign v3_1622710136_248 = 2'b00; 
   assign v3_1622710136_249 = v3_1622710136_62 ? v3_1622710136_289 : v3_1622710136_250;
   assign v3_1622710136_250 = v3_1622710136_251;
   assign v3_1622710136_251 = v3_1622710136_60 ? v3_1622710136_279 : v3_1622710136_252;
   assign v3_1622710136_252 = v3_1622710136_55 ? v3_1622710136_258 : v3_1622710136_253;
   assign v3_1622710136_253 = v3_1622710136_53 ? v3_1622710136_275 : v3_1622710136_254;
   assign v3_1622710136_254 = v3_1622710136_51 ? v3_1622710136_271 : v3_1622710136_255;
   assign v3_1622710136_255 = v3_1622710136_41 ? v3_1622710136_267 : v3_1622710136_256;
   assign v3_1622710136_256 = v3_1622710136_39 ? v3_1622710136_263 : v3_1622710136_257;
   assign v3_1622710136_257 = v3_1622710136_37 ? v3_1622710136_259 : v3_1622710136_258;
   assign v3_1622710136_258 = v3_1622710136_18;
   assign v3_1622710136_259 = v3_1622710136_36 ? v3_1622710136_262 : v3_1622710136_260;
   assign v3_1622710136_260 = v3_1622710136_261;
   assign v3_1622710136_261 = v3_1622710136_18 - v3_1622710136_38;
   assign v3_1622710136_262 = v3_1622710136_15;
   assign v3_1622710136_263 = v3_1622710136_105 ? v3_1622710136_264 : v3_1622710136_258;
   assign v3_1622710136_264 = v3_1622710136_104 ? v3_1622710136_258 : v3_1622710136_265;
   assign v3_1622710136_265 = v3_1622710136_266;
   assign v3_1622710136_266 = v3_1622710136_18 - v3_1622710136_106;
   assign v3_1622710136_267 = v3_1622710136_81 ? v3_1622710136_268 : v3_1622710136_258;
   assign v3_1622710136_268 = v3_1622710136_80 ? v3_1622710136_258 : v3_1622710136_269;
   assign v3_1622710136_269 = v3_1622710136_270;
   assign v3_1622710136_270 = v3_1622710136_18 - v3_1622710136_82;
   assign v3_1622710136_271 = v3_1622710136_49 ? v3_1622710136_272 : v3_1622710136_258;
   assign v3_1622710136_272 = v3_1622710136_48 ? v3_1622710136_258 : v3_1622710136_273;
   assign v3_1622710136_273 = v3_1622710136_274;
   assign v3_1622710136_274 = v3_1622710136_18 - v3_1622710136_50;
   assign v3_1622710136_275 = v3_1622710136_145 ? v3_1622710136_278 : v3_1622710136_276;
   assign v3_1622710136_276 = v3_1622710136_277;
   assign v3_1622710136_277 = v3_1622710136_15 - v3_1622710136_18;
   assign v3_1622710136_278 = v3_1622710136_15;
   assign v3_1622710136_279 = v3_1622710136_58 ? v3_1622710136_280 : v3_1622710136_258;
   assign v3_1622710136_280 = v3_1622710136_288 ? v3_1622710136_287 : v3_1622710136_281;
   assign v3_1622710136_281 = v3_1622710136_286 ? v3_1622710136_285 : v3_1622710136_282;
   assign v3_1622710136_282 = v3_1622710136_284 ? v3_1622710136_283 : v3_1622710136_204;
   assign v3_1622710136_283 = 8'b00010110; 
   assign v3_1622710136_284 = itemTypeIn == v3_1622710136_234;
   assign v3_1622710136_285 = 8'b00001111; 
   assign v3_1622710136_286 = itemTypeIn == v3_1622710136_40;
   assign v3_1622710136_287 = 8'b00001000; 
   assign v3_1622710136_288 = itemTypeIn == v3_1622710136_42;
   assign v3_1622710136_289 = v3_1622710136_204;
   assign v3_1622710136_290 = 8'b00000000; 
   assign v3_1622710136_291 = v3_1622710136_62 ? v3_1622710136_323 : v3_1622710136_292;
   assign v3_1622710136_292 = v3_1622710136_293;
   assign v3_1622710136_293 = v3_1622710136_60 ? v3_1622710136_308 : v3_1622710136_294;
   assign v3_1622710136_294 = v3_1622710136_55 ? v3_1622710136_300 : v3_1622710136_295;
   assign v3_1622710136_295 = v3_1622710136_53 ? v3_1622710136_300 : v3_1622710136_296;
   assign v3_1622710136_296 = v3_1622710136_51 ? v3_1622710136_304 : v3_1622710136_297;
   assign v3_1622710136_297 = v3_1622710136_41 ? v3_1622710136_300 : v3_1622710136_298;
   assign v3_1622710136_298 = v3_1622710136_39 ? v3_1622710136_300 : v3_1622710136_299;
   assign v3_1622710136_299 = v3_1622710136_37 ? v3_1622710136_301 : v3_1622710136_300;
   assign v3_1622710136_300 = v3_1622710136_19;
   assign v3_1622710136_301 = v3_1622710136_36 ? v3_1622710136_302 : v3_1622710136_300;
   assign v3_1622710136_302 = v3_1622710136_303;
   assign v3_1622710136_303 = v3_1622710136_19 + v3_1622710136_8;
   assign v3_1622710136_304 = v3_1622710136_49 ? v3_1622710136_305 : v3_1622710136_300;
   assign v3_1622710136_305 = v3_1622710136_48 ? v3_1622710136_300 : v3_1622710136_306;
   assign v3_1622710136_306 = v3_1622710136_307;
   assign v3_1622710136_307 = v3_1622710136_19 - v3_1622710136_46;
   assign v3_1622710136_308 = v3_1622710136_58 ? v3_1622710136_309 : v3_1622710136_300;
   assign v3_1622710136_309 = v3_1622710136_315 ? v3_1622710136_314 : v3_1622710136_310;
   assign v3_1622710136_310 = v3_1622710136_313;
   assign v3_1622710136_311 = v3_1622710136_312;
   assign v3_1622710136_312 = {v3_1622710136_217, coinInNTD_50};
   assign v3_1622710136_313 = v3_1622710136_19 + v3_1622710136_311;
   assign v3_1622710136_314 = 3'b111; 
   assign v3_1622710136_315 = v3_1622710136_316 >= v3_1622710136_322;
   assign v3_1622710136_316 = v3_1622710136_321;
   assign v3_1622710136_317 = v3_1622710136_318;
   assign v3_1622710136_318 = {v3_1622710136_217, v3_1622710136_19};
   assign v3_1622710136_319 = v3_1622710136_320;
   assign v3_1622710136_320 = {v3_1622710136_52, coinInNTD_50};
   assign v3_1622710136_321 = v3_1622710136_317 + v3_1622710136_319;
   assign v3_1622710136_322 = 4'b0111; 
   assign v3_1622710136_323 = v3_1622710136_324;
   assign v3_1622710136_324 = 3'b010; 
   assign v3_1622710136_325 = 3'b000; 
   assign v3_1622710136_326 = v3_1622710136_62 ? v3_1622710136_356 : v3_1622710136_327;
   assign v3_1622710136_327 = v3_1622710136_328;
   assign v3_1622710136_328 = v3_1622710136_60 ? v3_1622710136_343 : v3_1622710136_329;
   assign v3_1622710136_329 = v3_1622710136_55 ? v3_1622710136_335 : v3_1622710136_330;
   assign v3_1622710136_330 = v3_1622710136_53 ? v3_1622710136_335 : v3_1622710136_331;
   assign v3_1622710136_331 = v3_1622710136_51 ? v3_1622710136_335 : v3_1622710136_332;
   assign v3_1622710136_332 = v3_1622710136_41 ? v3_1622710136_339 : v3_1622710136_333;
   assign v3_1622710136_333 = v3_1622710136_39 ? v3_1622710136_335 : v3_1622710136_334;
   assign v3_1622710136_334 = v3_1622710136_37 ? v3_1622710136_336 : v3_1622710136_335;
   assign v3_1622710136_335 = v3_1622710136_20;
   assign v3_1622710136_336 = v3_1622710136_36 ? v3_1622710136_337 : v3_1622710136_335;
   assign v3_1622710136_337 = v3_1622710136_338;
   assign v3_1622710136_338 = v3_1622710136_20 + v3_1622710136_9;
   assign v3_1622710136_339 = v3_1622710136_81 ? v3_1622710136_340 : v3_1622710136_335;
   assign v3_1622710136_340 = v3_1622710136_80 ? v3_1622710136_335 : v3_1622710136_341;
   assign v3_1622710136_341 = v3_1622710136_342;
   assign v3_1622710136_342 = v3_1622710136_20 - v3_1622710136_46;
   assign v3_1622710136_343 = v3_1622710136_58 ? v3_1622710136_344 : v3_1622710136_335;
   assign v3_1622710136_344 = v3_1622710136_349 ? v3_1622710136_314 : v3_1622710136_345;
   assign v3_1622710136_345 = v3_1622710136_348;
   assign v3_1622710136_346 = v3_1622710136_347;
   assign v3_1622710136_347 = {v3_1622710136_217, coinInNTD_10};
   assign v3_1622710136_348 = v3_1622710136_20 + v3_1622710136_346;
   assign v3_1622710136_349 = v3_1622710136_350 >= v3_1622710136_322;
   assign v3_1622710136_350 = v3_1622710136_355;
   assign v3_1622710136_351 = v3_1622710136_352;
   assign v3_1622710136_352 = {v3_1622710136_217, v3_1622710136_20};
   assign v3_1622710136_353 = v3_1622710136_354;
   assign v3_1622710136_354 = {v3_1622710136_52, coinInNTD_10};
   assign v3_1622710136_355 = v3_1622710136_351 + v3_1622710136_353;
   assign v3_1622710136_356 = v3_1622710136_324;
   assign v3_1622710136_357 = 3'b000; 
   assign v3_1622710136_358 = v3_1622710136_62 ? v3_1622710136_386 : v3_1622710136_359;
   assign v3_1622710136_359 = v3_1622710136_360;
   assign v3_1622710136_360 = v3_1622710136_60 ? v3_1622710136_373 : v3_1622710136_361;
   assign v3_1622710136_361 = v3_1622710136_55 ? v3_1622710136_367 : v3_1622710136_362;
   assign v3_1622710136_362 = v3_1622710136_53 ? v3_1622710136_367 : v3_1622710136_363;
   assign v3_1622710136_363 = v3_1622710136_51 ? v3_1622710136_367 : v3_1622710136_364;
   assign v3_1622710136_364 = v3_1622710136_41 ? v3_1622710136_367 : v3_1622710136_365;
   assign v3_1622710136_365 = v3_1622710136_39 ? v3_1622710136_367 : v3_1622710136_366;
   assign v3_1622710136_366 = v3_1622710136_37 ? v3_1622710136_368 : v3_1622710136_367;
   assign v3_1622710136_367 = v3_1622710136_21;
   assign v3_1622710136_368 = v3_1622710136_36 ? v3_1622710136_371 : v3_1622710136_369;
   assign v3_1622710136_369 = v3_1622710136_370;
   assign v3_1622710136_370 = v3_1622710136_21 - v3_1622710136_46;
   assign v3_1622710136_371 = v3_1622710136_372;
   assign v3_1622710136_372 = v3_1622710136_21 + v3_1622710136_11;
   assign v3_1622710136_373 = v3_1622710136_58 ? v3_1622710136_374 : v3_1622710136_367;
   assign v3_1622710136_374 = v3_1622710136_379 ? v3_1622710136_314 : v3_1622710136_375;
   assign v3_1622710136_375 = v3_1622710136_378;
   assign v3_1622710136_376 = v3_1622710136_377;
   assign v3_1622710136_377 = {v3_1622710136_217, coinInNTD_1};
   assign v3_1622710136_378 = v3_1622710136_21 + v3_1622710136_376;
   assign v3_1622710136_379 = v3_1622710136_380 >= v3_1622710136_322;
   assign v3_1622710136_380 = v3_1622710136_385;
   assign v3_1622710136_381 = v3_1622710136_382;
   assign v3_1622710136_382 = {v3_1622710136_217, v3_1622710136_21};
   assign v3_1622710136_383 = v3_1622710136_384;
   assign v3_1622710136_384 = {v3_1622710136_52, coinInNTD_1};
   assign v3_1622710136_385 = v3_1622710136_381 + v3_1622710136_383;
   assign v3_1622710136_386 = v3_1622710136_324;
   assign v3_1622710136_387 = 3'b000; 
   assign v3_1622710136_388 = v3_1622710136_62 ? v3_1622710136_418 : v3_1622710136_389;
   assign v3_1622710136_389 = v3_1622710136_390;
   assign v3_1622710136_390 = v3_1622710136_60 ? v3_1622710136_405 : v3_1622710136_391;
   assign v3_1622710136_391 = v3_1622710136_55 ? v3_1622710136_397 : v3_1622710136_392;
   assign v3_1622710136_392 = v3_1622710136_53 ? v3_1622710136_397 : v3_1622710136_393;
   assign v3_1622710136_393 = v3_1622710136_51 ? v3_1622710136_397 : v3_1622710136_394;
   assign v3_1622710136_394 = v3_1622710136_41 ? v3_1622710136_397 : v3_1622710136_395;
   assign v3_1622710136_395 = v3_1622710136_39 ? v3_1622710136_401 : v3_1622710136_396;
   assign v3_1622710136_396 = v3_1622710136_37 ? v3_1622710136_398 : v3_1622710136_397;
   assign v3_1622710136_397 = v3_1622710136_22;
   assign v3_1622710136_398 = v3_1622710136_36 ? v3_1622710136_399 : v3_1622710136_397;
   assign v3_1622710136_399 = v3_1622710136_400;
   assign v3_1622710136_400 = v3_1622710136_22 + v3_1622710136_10;
   assign v3_1622710136_401 = v3_1622710136_105 ? v3_1622710136_402 : v3_1622710136_397;
   assign v3_1622710136_402 = v3_1622710136_104 ? v3_1622710136_397 : v3_1622710136_403;
   assign v3_1622710136_403 = v3_1622710136_404;
   assign v3_1622710136_404 = v3_1622710136_22 - v3_1622710136_46;
   assign v3_1622710136_405 = v3_1622710136_58 ? v3_1622710136_406 : v3_1622710136_397;
   assign v3_1622710136_406 = v3_1622710136_411 ? v3_1622710136_314 : v3_1622710136_407;
   assign v3_1622710136_407 = v3_1622710136_410;
   assign v3_1622710136_408 = v3_1622710136_409;
   assign v3_1622710136_409 = {v3_1622710136_217, coinInNTD_5};
   assign v3_1622710136_410 = v3_1622710136_22 + v3_1622710136_408;
   assign v3_1622710136_411 = v3_1622710136_412 >= v3_1622710136_322;
   assign v3_1622710136_412 = v3_1622710136_417;
   assign v3_1622710136_413 = v3_1622710136_414;
   assign v3_1622710136_414 = {v3_1622710136_217, v3_1622710136_22};
   assign v3_1622710136_415 = v3_1622710136_416;
   assign v3_1622710136_416 = {v3_1622710136_52, coinInNTD_5};
   assign v3_1622710136_417 = v3_1622710136_413 + v3_1622710136_415;
   assign v3_1622710136_418 = v3_1622710136_324;
   assign v3_1622710136_419 = 3'b000; 
   assign v3_1622710136_420 = v3_1622710136_451;
   assign v3_1622710136_421 = v3_1622710136_425;
   assign v3_1622710136_422 = v3_1622710136_423;
   assign v3_1622710136_423 = v3_1622710136_14 & v3_1622710136_55;
   assign v3_1622710136_424 = v3_1622710136_12 == v3_1622710136_52;
   assign v3_1622710136_425 = v3_1622710136_422 & v3_1622710136_424;
   assign v3_1622710136_426 = ~v3_1622710136_427;
   assign v3_1622710136_427 = v3_1622710136_428 == v3_1622710136_15;
   assign v3_1622710136_428 = v3_1622710136_450;
   assign v3_1622710136_429 = v3_1622710136_445;
   assign v3_1622710136_430 = v3_1622710136_440;
   assign v3_1622710136_431 = v3_1622710136_435;
   assign v3_1622710136_432 = v3_1622710136_434;
   assign v3_1622710136_433 = 5'b00000; 
   assign v3_1622710136_434 = {v3_1622710136_433, v3_1622710136_8};
   assign v3_1622710136_435 = v3_1622710136_50 * v3_1622710136_432;
   assign v3_1622710136_436 = v3_1622710136_439;
   assign v3_1622710136_437 = v3_1622710136_438;
   assign v3_1622710136_438 = {v3_1622710136_433, v3_1622710136_9};
   assign v3_1622710136_439 = v3_1622710136_82 * v3_1622710136_437;
   assign v3_1622710136_440 = v3_1622710136_431 + v3_1622710136_436;
   assign v3_1622710136_441 = v3_1622710136_444;
   assign v3_1622710136_442 = v3_1622710136_443;
   assign v3_1622710136_443 = {v3_1622710136_433, v3_1622710136_10};
   assign v3_1622710136_444 = v3_1622710136_106 * v3_1622710136_442;
   assign v3_1622710136_445 = v3_1622710136_430 + v3_1622710136_441;
   assign v3_1622710136_446 = v3_1622710136_449;
   assign v3_1622710136_447 = v3_1622710136_448;
   assign v3_1622710136_448 = {v3_1622710136_433, v3_1622710136_11};
   assign v3_1622710136_449 = v3_1622710136_38 * v3_1622710136_447;
   assign v3_1622710136_450 = v3_1622710136_429 + v3_1622710136_446;
   assign v3_1622710136_451 = v3_1622710136_421 & v3_1622710136_426;

   // Output Net Assignments
   assign p = v3_1622710136_420;
   assign coinOutNTD_50 = v3_1622710136_8;
   assign coinOutNTD_10 = v3_1622710136_9;
   assign coinOutNTD_5 = v3_1622710136_10;
   assign coinOutNTD_1 = v3_1622710136_11;
   assign itemTypeOut = v3_1622710136_12;
   assign serviceTypeOut = v3_1622710136_13;

   // Non-blocking Assignments
   always @ (posedge clk) begin
      v3_1622710136_8 <= v3_1622710136_23;
      v3_1622710136_9 <= v3_1622710136_64;
      v3_1622710136_10 <= v3_1622710136_88;
      v3_1622710136_11 <= v3_1622710136_112;
      v3_1622710136_12 <= v3_1622710136_131;
      v3_1622710136_13 <= v3_1622710136_152;
      v3_1622710136_14 <= v3_1622710136_170;
      v3_1622710136_15 <= v3_1622710136_175;
      v3_1622710136_16 <= v3_1622710136_206;
      v3_1622710136_17 <= v3_1622710136_220;
      v3_1622710136_18 <= v3_1622710136_249;
      v3_1622710136_19 <= v3_1622710136_291;
      v3_1622710136_20 <= v3_1622710136_326;
      v3_1622710136_21 <= v3_1622710136_358;
      v3_1622710136_22 <= v3_1622710136_388;
   end
endmodule
